��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�C��vU���Z�
ɠI�6t�s$2�@�c�5��v0���Vd(*(��O�(km=`���/�H��$�s/7F�6+���לE��f�r*��1�CֳEth�5h�P�w�7�ny'nJ<���"2nߴT���B���SE�>VL'����3H�DJo�Jʸ��O}_^�% }q�����\,z��rg���;gs��~���"��I]o�*��0J������r�@�7�'����?��@r�6=Y^{�&h*x|p��C=���fq�Wkڐ��p����͠��M{8��p�����ҋ�	����o<f�ю ��:V��i���$�\.��|�S�!�Oj��*|�T��<x���tZ�ǀ6�B��L�I�#��TX��N�M��?1�ci���9����,�s`��5����d
;�V�G�LZ�R�F-q%�sર{�cI��ѓi��$2�@yF��2w4��P��*G葐��T����Qg��u��S����)b���wl�ڶ�4F։�Y*�j������]��)8�͜�/~s�����	��r�Ǽ��A����`*d���W:H�:,�4�ṖE��A�����	�My����j��^/1�*x�ar����j�$���ڷ]��'����88*�z���������	utpDѫ�y��� m��4po?�)��&w�X�x����V)��C)�y����
��̱+:��*'�ix��L�N����H���(����X��+�hXD�*դ��Q��n�,|��lXt�wF�r��'���p�1�C&�~����Za��)�d!��FvJ]E� ��*�}x%�ܠZ#��V���<c�Q��\A���,���^�哧z˴j��>�����A�s��u�&4�Yo�b�'�#8���?-��B=��*������ʿ��r�bc���)']�lV�E>�a��9�a�P�k(t��׎���gil�u�[�ŉQ\(@Ư��y�<��<k����q7)�@���8UH����	��������B�Q��y.�F���lS��5���>�&%֏�@@5w�᫧;��.��R��.��G�5�C:�Io3)L�|u��������㾺�bwtIf����)�UӝОvշ��	&��>(o`NҢX^��->���z��V��q��jӅ,j��"=�y�F^H�&�m}	B�ڐ��>@�<�Re'�F�8�͗�� �k֝z��a�� �q��?���r
�?�q`,�N�=o�7�z��8<g��>������T��=���^��F%:c���S�h�r��q
P��]���#�-O��/�T��.ָ�H��\{�V�ȥ���);��~����܉��0~0�Q�K�B�n;B��+��'x<��s��і7��X%�4򑡘
�W�=�U?�:3ŽXi�yu��[��d���k�B1�;��ޏ%�FӶ�hn�݀;J�7,"V�J� �m�L�G��*�=cbݵ�h��Gvԑ���צ;��j��\<})�h�� �zL_4d'@+1(xB�$L��9YR����D�"�c'6��͏T�y�U%�NTA����A++[�W�/��R���R�}� xZ�f�6OQΕ�k��"�t��@���S����ϸT��22�TO��� �A�U�A5u�C2���r�.���*��oZ���}](�QE���EJCæ*3��#!['h^Ӕe�xS'��Y�jQP�	n�����@�1�o�e���j��IJ/y-�-"�P�X�攦w�D�^?�R�T��|��I%]�v��PxáΕ��h�DAZ36��MZ!�@C�n�ө�\4��S����گa��a곿����������(y�1�^��⓵���w`uy�����"��6��w�����q�>g�ĸ>ٮX˜�S/��/u��^�΀(��`fM�>�-a�y�J����r��j��� �4�sk��H=Xk�@��K8�^���"��4�	�x9��_|	�IN�?�B��Da�6y��܌n�Q��	H AĶ��)�MƆ��B'$ �*���C���|Z�����QE(-��[��/,Gmٮ*T�݂��F�>
���2'"�rk�����t�C.*湛h��\�v�1�F;��esp����]��i�@�ՙ�o�yᙼ�����0Q	�]?�5� 6�(�8��K�ph|�ᙆm&ŮF�80Ұ53
O�i�*h&�y_~�G����I�T�c�4�X��������v5}��O+Ҷ��y����Rv����m���w<��T�hL-5��
03�jv��0q��G"�a)~��{���j1�w `�; 3������i`X�%���?����@�#�^i9D�bw��1���<0Ɍ ;�lUmp�� FƱ$�x�U^f�B���Vi�n�����{#]>8C^�VSp�$�>1qb�3^9P�	��?a��g����I�HJ0�?���o�����i(�Qh���r7$	��'��~2�d+{q�DG�
�1�%p��.�w˷P��,"YZ� �Wg�(��]Jn�g��䛋"uu��,�qR��;o���;�X�����/��-[��޽�j�t���7�K�I��s��a�<��f4�D.yx��|�PK��]�e�D�浏g�r��;�Pķ�z�:��q�Ϡ���8D�����U�5ݞtn����/�э����.{�'!�]<2���96�E�h(Ȕ;&Ծ?���������t��W[�E�K�x
����Q �U1F(2V_k�^4n��u�˿�z#6�d`��T��H�����c�����D��݉z�r�SK��)���܂>����V�F_H��P��5��j����u���!&��wQ+SD)���pO�/g���<��۟����)������R��o���ET����.��Z1XI��ǐ$�Z���%���/��� �5]�K��[;������G�`�t������vfjty��B:���:���+�(�5H'���;���f.��o>��a�>:�]7+�0T`�a����qd:d/;%�@�j <bs/^�C�����PN����1P�B}7A0�U����ی�b([h]@������j�	���d�S��v����mx����H��9���L����]�t�ԕ����E��;7\�z��"\����	��r�K��0V�;���f"�s�������(��]uY�;ŮH�����>@V�u挌��I�WK�$���n�8�Ť�1	���ZK�/����l$��-@��>����
����>vS+j�@>��A���Z��g�OM.���W���5��8�G9gb�p��SwE���{�m�n��C�_�6�l*F��/�r�5M��x�Ԝ���egkc�4���<�'f*_p�T��ÿ8�e��n�Oԟ[B���A�>u�S<�)lZ��3��,Sv�T���H�:��g=�SC�ߏﯠ��Z}j�(�ϐihNWa�߅��"3PH#՗�c֊�p:���ڇ�lfPya!���3g�VJQdߍ"�a47�U�J�*	���MT��@��X�g����Wx�ξ�G��fi5�e�oTܺ�n�8��+괸�g���&��%e�MM.�7��
r��Pw_�.Zr���
���Oj��P)�*��	������Փ!��F�~�S��ԣ��F����`��{X��pѠ�Hg}��x�Mol\�~R�6/�"d��
���I�6�n,�Wڙ�$i$�vs�}ݛ% � ��-S�f�~�AZ�N<�Q�#t�:8�1���Rb}�'�OxN����̚^J0����W6'� ��mo�`-�|�P�_�[���K6�����]*$o��ǖk�jt}��W�^1F����M��b��C���x2�_�b�~�8 �����2q��y�k�E�U�I��UMn�6�Ɲ��]��8D��	o��uT��P���MN�e�N�]�ФL֧���>{��OLuo]���3�֕0�_�����??����8m��@��R��"K��C��iFT�ꦯ���Ș2�*6�	/&� E�D��gIPv���v�+I"��L�Xd���+�����*f'�".]����\k�@m�H����S�?�j����G�h�~���˒�������
�P��sӵ�<��
�PS�EF$�w6A��/���Ί(Q
y��c�S6�c�j�������G�}�\w3H�l�x��Ks�`�Go���ԩ3�B(k/�I��U�]_�C΂&�~�`>>�P��2�<DnL�"'!�C9;�n�'�)=�O[( ����6����t��"�D�jQ:���r���	��.��V�p����2��E�W��-ð NT(�رI0;%���
0i�6|��\9���k˼�Z;H{{��,S^qI�����?=̆5@�E�_	yFp���QK��Y�����{��W�m��U��:U@�B�
�L�ˠ%Rs,�=һ1/� W���l������=�5 =���Vy��L�d�}�r�V �_��S�䋐��"��cOY�����C�%����_�Ã@��&��۰c� �7\:q1���~��fÉH��K����+�)4���3�)�oH�'8Q"!��_�u��P�lr�'��e`��f���=Ua5-�(���=Ɂ��._��P �wfXzC�m���W��XH��_��(����8J��2┘�nUUt�HR�gk���Y�#�=������F��]ĳ3�%��y;������ar�6#3�Ȝ�r����A\��A��`ʇ�T��ѷ94�AX��` 1���� ��^F@=ם�lh� ��F����*y�؉`���Y�I��}��d^{�w�ĳ��+�����׭�s�9�e2O�#��@�:'��뽎gr�C�eWXҲR{;@�h�ܒ���Z��b;#	��W갭a����<��d �T�Ig�e��z 
��n:�$�3�\	m�个]�I�?��-�F�0j��I2���W=&�W3�؞���.k̭���q��]A��p�q���p
�y��r�S�C]�� �1���<��N�@R�`S໳/|�ӆc�!@ba��L	 b��.M6X;P�C.sUxT���؂Y#w�TcR�2ژ�,�fuKll5��Y�kD��@������ж+�PU��������#�I�[�������	F������r`5���+{d��t���h=ڏ=y�t XE�+.�^v2Ĭ��l��b��F �*�K��N�J��cn	i�3�z 3������qW��E�@M�Z$b�������{U.���hpB���xwd�#���N+�4�- ��߽� �Z�l�W��1������@���`�np��t��!��H�Zg��/h#�|K;�$hi�PH���ӓ��	����{�'vrP@�>ß�,W!g�G(�2��K�u5���F��se�$��{?��<�3�[ �z-a�t^Od��qiؼ�B��`P���D��� ���$
L%7E>^WJ�ٔҡ�*,a�+4"��C�-u9ER*����"�Pjߋ�F�Ƃ�fX������lR� ,ܦ�v���ԯn��eD� ���6T?Un|b;*��s�=^k�0E��7�X���DN��}�0��w�� �U�.���˕�,��4��6�-��B��?qw6�����dO?S	}�׺�`f���L��to��]G���!��F�F�Tn.��aJ�S:,j����Vx�	,!q4��i�����fr%-��*�� �ڲ9��w�I\y���Z�l���m�O��f�M�!@Zb�*�9���[8����L�@����A3��d2�%@��=t��� rJ29 �k�H�K��J�qC�ѨŚ��@ͳ(��������2���* ���8�x�1@?D¨c���N��Ļ�?�T��^�c
�&�U�^ãW��d$N�a\����5Y1��ʚ�ּ"Ɔ ��Ȉ���x7v�VI5Y���0'���&}�^LE��8�$��b�'f�m'�'���h���s}+}��ϳ�7�]^-���t��Ɵ��@���"CM����}������qL=�b5v�ÔJ&��d�Qԑ�_Q���OϿs�1�I��PǾY��!]L�u_���1x��iA����*�>t���\ �jP���
VB~3��GJ�_�N�Q��P�лC�Ѫ*3��o��bw�������ȋfK��j���6��~�®,4,��:׋帒�H��c�O<}���H��腊ׅ莰���`����G>���":<|��Xe�*�R-ݱ�� v����O$"�o�c��B���O$�e���A����E0���z���k`K���Í�3�*PB���J<d�B���RE�y�B}�����⵬&�k�e5x�;�7�@m�������qYI~��(�(���EM�NjJ���9b?A������:���L�TTRH��T�>]� `�� �xI�[�P�8[i���g��Yc���X�2�\Vx*c�9�(7�X��
��(E[�3�PT��'��|�YW��a���h��v����Ws���
�~���y>�u�Jy�x��IW��`K�,��|�٨�`+��@�N�x���feBo!���߭]���ǂ���T�C��yl��O�)���1��#�4�P�!(��e�(�M����,���5v�o4�sڒ�)�)����̷A���4�e�cE��'�,R�
f�n����q�3��L����z��17=%=%�z!�햎`du��L��u��8��lG*��@pph��Vp�;��;��ib�~1�y�
���.t](:LS�ɮDxf��s^\&u~Au�^����b�AI郛x�{���L\�X�V3 �V�����aXX;�6o�(\G��`��Z�yn��Exg(�al�(s�2=�}آ�{��3���W��b�f/�J���F�cW���HU�Χ/~�~���ŝ�Z1Ĥb�����3����*�a�l��p���"���� q���D��7!V`m9�\A�H;�}�����6��`��߄��i{?�ݜSw6�rU9Tp	��$�~?��d���ɼ�O<�2c����	Б�P����;Uޛ�F�e��7��*w�OR-I����W$��%p��;Ћz���o�!�B8)
e��F��x�Y٫����#��!mL�<{
�I�X%E�w��v��3��;�D7�T�9�e�ZK�O�h���� ��<�;��pJ�s�����Z�Z�ܸ��AC�,M��\���W}r	��8U�@	g �ڪ���yr:�X4A;��ݣâ�k�<��}2��/��(�B�����0t��rr�q�'�)24�ׄy�#�s8�O��B� �C��]h���99�� �Ie������D��v9�֑��P<� z5�����i�;S�x&?� 'o�=	V� /����e�TOSL7�k���}�^k���Gr�
��)WQ�&�����q�EEm�����	Zؚ.�� �����=&�bp���GL���=�Δ�ഖ������������7�&��Vֲ5��s�_G2G3�&[oa���[��ҳ%N�Թ�w����%��t�S���E����z��T��
�4GaȲ6Y��x��=���aT�q�M�*��j]���J&��<o4�s"��=���EH7t�ѷ���d�{�ʼFӞ���P�x��a�)�wɚ���[�N�)X�׌��u�3�%��_P���z�\F�=&k����]y�b���k�J�I�mM�@[�IeO�=}znQ2V^�����=��D�%;�n��7�~6���֤.��D�Q��Oŗ;�g�wY�T��53��{7vk�`�3T�%��yp7͛#aR�E9SR�d�8d�a�.D2&����HЇ ����s%_K�xC�#~�'nW�/,��H/4��vѮCj��<w�y��M@_sY�~�����(g#'<�0�(��_�|
Pϣ$�bB,gUKߨ=�4�
������_@�����0��s������c��Y+C&=��Ғ2�7 Sw�"���<,-�"��)SU�4Y��h�z]~��Y/�������"�q`&߅�JhL�ӛ�/+�0�� (�k	!݆,�F����A�Δb��rt��	����ag0��Ya%|��@�۹}�Έ*�k��Q�cƦ�n@�P��9�����|E҉\X�}�J�tj�����iL`��~����8|�[s���L��K��v�W����m��p(��NWn���}9����������h�� �TK�����8�0�<��~���� �#������>�B@V��r��$ڑ�Ph��'�)��@��Ӊ�4fwy�?j{-O@��<|���Ĵ�%cI���Hm�Y%�=$A(x��R^��f���
��E�*�]x+�*������5��wN���/�q?0v�"��F�g�Ll݂�3�h�Y��Vw��=Y�i?h>P[ܻ.t�u+NG�z*uwG�%�T����3���{�\�� ��_=o��,5����=�8�D��cG-���S��Z�G���gn���M�dɝTA>b!�*-�3p��a�#^/��x相4�X�~�=��&)߿ �q����&�Ag����wވfl��K����n�H$/�
,��+�a90��P���Z9���݀4I �k��<��-���� Zɝ��B�ɾ��UF�4)�f���HC��5�l����,f��Ѕ5`8E�C��)����<�]�P}`�R��������ZT��lw��v�;�1sϴ��֟���a,|�wʅ�:�vQ����� �Iv?���/O���դ>v������+=� �9kKz0�4�7'����GP��l,,&{�6;�É�����D���L�W����B�@N��m*t�F��C]�Hu�.�P���x�cO�HTiY����9�{��q�=F숹��v�Q���b"~��Ugi�.2�Y(�%�:e�f��'yη42�
z��V�e�
��Et~s#*Sj̽�wyCD��,��l��.%)���[�Slo�,�����E%-�Yx8�]�1�ɰf�܋";'�|.��;�ƥ�����Q��7V����V�����t���G4�\�z�X��x��قT��w���t�2SYN��ݯ�g�i��	b،�^{���UJI�iD��W��D������>� �kf����\1{ ���z�ήro
۾N�M�uĞ����s��T]�LK��K���RT֘N��C�o{�e��`g��Zɱ=5��$άIГIu��/��
' N�|	��A�w�8��
X^{�N�t��	��{�:L�W��=�J���7(�$���ڈtC��ڀ�ΜN%�ie�0㱜;�궠����+Q�Sd�]���AH��
��X��#"�΋��s���������z�����o�d'>�r�Ĳ�V��l=���̻N������ơrc?R�T��I��g�v-C����bn��K@�[��F�K���W���g7j�����)\jZ;���V&�/lt@���nlI]��uW$�s=��K����Մɣ[Ap8=]������=$��)��k�KSf�"o�>�������ܸ�������TJl��.%'�W��a�	�g�0;��)8]=JM;�A��KD ��4���^l!���%wSG��}�� M�Q��U�6��[h!|�#`�5L��kD�ӥW�Τ��%�9]�L��P�ją]E9�k����3�2���ّRi�=���Z�F���� ߚ�Px7a	V]��Ӫ���������9�z�S%��y!��b�2�YL���\6=���`�V3 �]�E�l��o����l�(aDvh)=,Xx��s�[�0毾���&��`x��|el�� ���ږ�3JYQ�q�B���_Sg�5ُ���Lf�.�#Pes_��X��E��
�ezj�XB�lg��:�!�(�`����=Y��~�V�s͋G�� ���囟tV���b��mC~d���Y�_0<��#�+8Zo fMk�S1�
���6b7=���(JD]�.�k�|���q�& nLQ����Z��N�-C謭m� ȥ��eM�c��
og{����,נ��/dՑ��o��f�����[O�؎�}��Z"|�;���ܛ�)���ڏ8�Yy�:U>l�Q�����w�h����cP;�����R"�E����D��<[R^���b���9xpg��3W��H?��
���x�z�& �M�[q]�=YT�0���'l�����y1��U�-�/�����1�$�/%}�"-�М� ����j�Q���g�C��Z bz���%����"�����:����~���gP���u�8�5z8b�T;g��~f��\��Eic-2eb����������s��5UlE�5�˼ z��#
���z8�E����32f�,p�4f��I;ru��	���A�~D�'�q�J¹Q/�`I�Ae��nuz�P���f	�a���z0�w�F���@��:��Oʛ;��_�_gEQv��Jd(�YX��'��e�B�[WL�n��8����lszj #_`T�
��H�քu����cZz�$4/.%�Z'�8�*�0�Zg�B:oj�Ggdz��9�HN��a)��� �<_y��`�ӆ7z�E=��"Qx�O��=[uiL�+�P��})M0+hG�8�ve���w�>���D*{���g�bSg�ۏ1���+Qj(��=�t75�H.c���Q�����}���F�z���5z!��	�ۂ�k@�������V�ZbUI�QL�Z�a�P�8��2
`5Rv�Ȱ���5�A!찺`���"�Z�#�O�R���4WR0R��<�Η|����ျ���~B��;��ו�s��;�w,Q����!�R9�� 1x�	���g=��f���jJĳ��� �< Tz����e���#�m���Wg��B��W�d_��)nhl�|�����tzNʜ��%��D�{ \�X;&o��3C*y��wi9�i�(ߕd� Xv�N�kJ��W�b�!�x��EYs$�O�q��řny'� �V�Ьh�S����!d��׈�[��!ˣ��5j����
� rV�/7�����kjL�@�z�����M2�A��K��