��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>Q�y�`�}����ż9�_)����������ꩪn�||��}�}9\㌨.���tR�±��R���ۓ>Wb��E#��Y&F��:�m3��Ybz�[��x�l�1èd@((��F�
bi�����V :���E���?���U�,�IF�f�
I���,ݴ3��91��O����"h�Jn7��G����m�Q�<IPWx��N�3��.M\�0?���{Q�h�pM�$I�薵	U����O-ʃ�։��T�p�y���Y|OZD�@;ꕰ����9�>"�,�0C��]�1��*��p=n9�ح`r}}Uј�i��!F&�_���񸷙@
�K[��%����׀�[u5
��À��EG&��k~��.Ug>D�.,P���]m�g�N��c��R=���a��V��b]� �+6m5�T��f�����nBc5�ṳl�[4��w�(�O�cMC�ډ�>�<�e���
ׇ��t������S��|�s�艨������i5|���^LC��� �,�����t��z���,��OC\�����M�;2tV㒋����i�K1��l<����ǫ�B�מ��+�p�Ɏ'�N���CM�{��-�������<{*"M����E����=^�w���`D������	,?���&-���#��D�o!y|��}��r��&��.�?.���u�=%F���/an��n���쳣B]�Qk�+�l����Dn�"��>�?L���(Nvm��	Z��!�:�u�C��Ԓ�Cn���0>�C�&d�W�W?Kr�f��.&��׎3����i��vn�C��Ea��9߸���o-��o=����+�a�8<�͐X��pp�[������Z��A�ǅZQ��;ys����]�����~�e�Ȥ���u����|�)�9;�ov����d��.��!)��n &���1����9��M2����ݯ�I�,Ada�P�L�*ÎgV�u�fY{M�ŭ�k��tp�t5v����r +��->3�E%()�u|��GW��o�f(����%}F;�$O\c�@��斡�kL���7�*�����ؐ&-dQ��,�a~�8 ?Z��5RqE	�� ���>_��QEF� �(��2���Ok��Y"o���V��m�y99�\K o]1�fI�����#9Q�a���K���d�b@u=�\/��{ �p�Z-��h���&\1v�G�)� k��B��zǢ�a���cs�q8��b����s�ѡ4�p3Z�߃�=/Ğ%���f��6����,�������Z^R�薶���@�*8��~��/>4d:�2�+p	���<v?] ?��狔���Ȟ�L|�&�i��)3�"֭��׊Mv��������Z-í/�k5�U��L�F���Dd�6�j�o`Jt@jvܣ۷�����Q;��T<D��ԭ��O����ϧ�w��!P��b]�^A}8N�Q�����f��P�dl���>�b��ENxZn5���A�+!���"���<f�*�/�$ã/`��O;�P��-�1�{�ˉ�$��8M���6`V��Dzɒ(q ���SO��nx+ۢ�Iv�zvۿ0���瀨�jTa��_�pU���2V���O\�\�._-o�W{9�KP��t��>���,��@��­V<�N�}�O܏�|6Bm<�RUcO���^J��/�J�"ļ�Ԩ���|��Db;>9����h����XR�Х֠�C�d�Eu���5WH�݌谯�O���?�f��.9*eP8(��A<g=D����ί� /��+�Y����� ��3Q���2
�|�/X-��
�YM��Y�{��2jҵF8�����\w%sH�?�-��_���Ǒ�e�;%��:
1%��A)9D��3�}�YUWہ8͆Ul*t͂�|-��G� #�g�r�����H{�������4g����p�Q^9e�: 3 ���l`�#^�蔌VP��u��#�/�ǷC;/�<��Y�g�e���&uF��0�A.��#��$^WO�5H��r��={��]y`�c�1���:YL�ւ|��'(2w��>�dK��I�*,TY��A��O�i5��Nn<7Dn�����G������
�{Z�m߰���C��r�="̓����7��P���?n�����w-����ۊԞP��=M�a��P�����D��A6Z#�s�Q��	��[Y��W�����6:���)���1��~9�F{b"��������(�뾗��`TKp>J�Ȭ���ZQZ�E��֗��?T����g��8(Y�&��W�(�V9�	_��T��i#���T�9��SJ����kzp��рIY��,k�Ȥ~�N�����������y �?	3vIN�ґ�'��U�7xG��Y�W�C6��G`ū���(�JӞ�e������W �������sO���f���싘ڣ�3'��D�ߵl�)8��7</Ջ��_Ex�nk]2�E.�5�;�3G�FS��J_#��!0�.��`��d4[^�j2�V���(���
5�㰇7�K���)x��X��oh�*D���A�)�3�Z����'0?z�v�%,Q��^j�q���
�s�Bt�D�Itr��X��Ľ��X��IC���I<3��y��_�Ʉ�W�i?��\�iR��J|b��ˢ�-�Ƌ��'�U*��l=��An(.9bv�u�ǆ�0ؓd��K��E)l���H�>��o~���� �dp1�2�lQ%�i��a�E8��F�rTy �!�����+1�|qOԪ��$���ӈ�X�e�m�4��9"?�l�ʧ�A�b�R�F�]�����}
���=�w��nb�C& ����:�
�<; ���26UE��e��O.V�3��a�K�њԱNhG��|������k����!(��t��GH���_M�X�hn\������2�(���[�~nǡ)Β Phn٦<rN<s.�͊$�W1E�1��Ob�zf��]�E����Aݤua�����̉���V/N���V7Q�/��{�篿�$ճʙ��k��續���*�Ϣ�!�[��(��* ��P{�D�Z���}���ڣ	ʂ`���t<�g��6{�sr�h8�Śxq��\�ݲ��7�9���4H��6��������0�~@�������pP.�+Aw���P��Y�'N獺1�\���HA��|$m5o�\����|WȎ�UZS�!��%ͯZXooԿ27�:�����s�v,�-т���ܕȀ�#�x^�͞�|~�>�K��h��e�R&��?߀��љ�Ȁ�T[�ocq&��N^��6pT�d�z'vJ	z�|��	�>?��m�_�Y�j�9�Ҷά���M��:Ql����é�SpI&��D�T�8$=�k�6�*l�H��ŀ�j{��m�A���cvv{{!T�Jel��dX�'�i%,�E^(�{`r�i� q�x*K�[��S!kNIM$�1���_��	����Yq�����v�3*�i���(�^���N��Z��~c��V�"8�>���o\�A<F�%����T��5j�rh=ʢz�������圓GHl�vM�T���y3��Dw��i��d����0�d�<Vo��[L�ܨ�T��رI }�B�������P�����_�e%�.��H�E�4���ȹ���O����U��끑b�T���X�2�v�<Y%��E5�F�@.Nƍp�T�#.�@��`��~2�G�v��U�{�e�3	�C�خ,����䳀����9i�gO-��!_�!UHpn��@B;4��0C$�*8:��o�]rp����0z.?���c�kg�8�`/U��"��( ��=;VХh��|
�I�4�:[[x[tْ%��#ڝC�*��݋�Dp, �,uy�9��@y=���.����s�m1$e;�Vh��������
�E<��Pg��1ad��'L����Sx��)���J"�1_�١���%(G&���@�*���;��Z�Z*���������?��"��Q����p>;�2�h�d�$�|*L
���qmOE�l��.��������L�S���O���P��08b��B�E'���\�"$�ɉ4]pJ~M3�*X��i6,J�_tQ ����퓦U|���L�t]��X]:ot`5������?r+��pD����y��N�M�JU-��7�E������E�w��p7�����Ȳ }��i^�cX�E�s�Fm�'I�
r�L<�@T)�ћJqM�kL"����t����j������6�i�H~
o�`��aσOq��H�Ƹ���TYK�᷃�h�v(!.3�d$ױ
�WV���O���*g��E��c}�J���K�땟���2$iR� J/����-7�s����ǅ
��4 Pѽ_�k3�+#�#>��>����GN�>��75�Dm��g�(CK���"���o�3d�up���7��B=6p8+�o2�o �Z�@�>b a���~����ЁAT"M��������A�Y�j*cB���W�Ze(��@c���NT�����@�%��ϝ�_#m�.�J� 㩙Ӛ�o|;���?� �<��n�S:��A��
0�Ix���P�]���͕>Kކ���4���S\��ߋ�竺��O�x���'�@+�� V�Ejt tK�^����no�|c3������0^5�K�#�C��0p8#�1L��qDUv��e�L,�(�ޛ.�7�4a�GĲd������^;�I����#����W�Z1�O����W��������uh6�E��+I�b����R�r�hY��z�����m���J(y[�!4������j�7�Ū	E����Kй�D�c+��S ن�0�>S���.h)�h=]7r=l�"�O_ε��X�OGf�UhI��u�`�VS4��k�)ƃBw��Ĕ^|����e�rY�ˤ��6N�[;��]͐2��|�1��:�㗿@t�勒���ﭔ��7)|VC���Y�ȼ�v'���Z�ܟ��<�����?��V�)�.rxZD-��y��x�tAS[�w3�$��w�o" Y��#Gߨ6=K��X�3�ulmlI~7�S]Ȼ��xZ"djB,�wj���t��x�/w^�hǢ�Ğ������̪�-��9w��#��8�����⮔���r��~��M��i3������s�1Qi�>�/�5���u��`>$|��@������G�W�x��C:�x�v��u�����袋���<���\��r]:���Nj|j��r���.eqOH¨�h�"����t�$�[/	V���\=P32�Zs� �^N�m%�ёU"�s׊���_�����(�^��M�/6p|gF������`���/+2H3���]��*�����K����P��p��zђ-v�/^8�a/Z�R9͋���1�J�_���G�JMK���cU�2E!�^#��W��-`��NBT7�r�C��$*��.� ����b�Sؿݺ��Țw=�ߜQ@1}c�	������/�J� x��LS�A��/o�ш�Q��>�C�����V+-L"4H�*Z��t9%�Q<����b?{�,#�*��Q��S��{��2ΐ�� ��N��[�_����'}5a�T�r*�q$��<�q���M���T<#á�z������	�Yx~v�������o���&����n*%3����R�+Q /��)d�*㬄Ihh�B"���#���M=ӎ
CA��.��,ڛ��7� )S���rΥ�����	�K.��+i7��7[� I��-	����Y)�_����'��o�B0@����@*}Ѝg�t��z�!i�L�B����
� ��<���q 
F��7�6ݟ�W���: �yp�w����o��^�VcɊ�4+3���D������)�楿Vm+g\�޷��N�$��X@��g;�jBC������¢����d�s��˻7�1��
�[u�5<�9D���昔���*7!x\{�:�
�N��J9r+4i�k�jAgg�֓��w~K^�i����Ռ%�#���겁��w��b�#b�V���w!s��B=�᳃7N/����gzS��օce�S{1ѺrM8�=�����4yC@�\�qYȈ�����sy�"�|��EjYOϙ����vآm�����RTu�.f��
�su��'�ī��J�;,HU�=2�ˉ���"l+(�%��P{rJAw��Oa�a��((���;"@"|9�M�K���6�^l�5��#��#��;�b8�ᳪ�E[JT�p�2�����a�d =[�|��u�9�50!<w|�^M�ͤ�P��j��\��F2rB5���=`�+���Z�"޼�bó�5�ɁuS�C���	��T��P�uu�G��2�k+�r[qЪ�s�*�|0,��Y��������!S}���80����hH�����D~&+�s�Ϟ��P\^�m著l�	]XUا���z��R�ɣ�v�gР.�����_̶���%D���6眼ml�9�#@�s����j8<\>�_�r���I�k�x�WK_��YP׽�Ľ�VdE�mc���4��� %S�iT˖))�,�_�O�,��o[QL��;��\��}�f�`܇S�a�fneZ�����z\(_�o`>�Kr89��!<�ѫ�d��{\o�g
u=��w�2CE��+A���=��+�����美*]�o'������wN����P��+�V�{|��:@�qS�����#y�厯��2�����'�h-&�
l�<iwߛ�����?|)�Ya(�2oɫ��C��E��=9YaDVđ+��ɮe�RY�%������A֊�U+�IA�]��ZO�ZϿ�F�1{�Ԧ�Q�~��H�x{>�]M�=Q�"������#Z@��AtUפ��Z��6��ɒZ~���K����%^�}ɗ�e�M����$�a�}0�[�u������� ���kX��J��X��&zl��!:��řA�kV��6�`��#�&+*%��W5U&���K�mR�	8k�X����˔=Cfe>�۠IgA��Xsi�5��f�@��;�;'�9���3�����`/C���y�	� �k��ʾ�*��~F�3����S"�<�"�x�h�@5��#kAnk�d���ENA(���5����-�p��d9����,�m+���l�'g�����j��/I4b�DV���1�>V�s��/
Y$]K�|u�y� 85i��*nx�0>aE��Vp���g3~s��ʸ]�T=�|`9�9����r�i���$$�X,`QL�^����}$�bW
�d��N�y�A�S�r�.g[�l���o�C��?���:\�mnGo���L�-��B��*ٔCB��`�Yˑ�"nEu/��k|>���4������5T�?�x�ݶ{�!�)֋�DnJ5��#

u�J��c�ݸf��i�a([A�D�N��IF5��9��i����mt��2)K��v�`,3��O��[�~=�V�]��$OT���&��,�a���E���Z�|m���C�����8���v% �3�k�دQ,��#7�?((�l�xe�!5�wQ�RSL��')�-G���OK"1��g��5��i�ט@����U�<X$-��m+�"1(�Tc<`��0�ߍ�	/H�V��,Rz���u+��P�\�ځ��f��rТ�+�>�bW���x��u�j�;t��Ϻ��Q�c`�������T#��3��sn���ݣn��R����b�Au*LA SDfRZ����70��9�C�H5��}�u5M�����`K&�R�6_,���S�.�D�X���!���Т�k6��O��Y}��M���x�  ^-�8��x+���`�c��Ǟ+$[0T��dY���ڍ"�f�E2(��9#��l��B�tѕ#UN��}`)Ǡ��ԗ��Rt�_ ��n�׊M�k7Aa:@��C�Er�#��
Z���9�=
ب�Vxz�z?�|��O�X�ww�V��Ҭl�?*^Gxc�ݘ*.B�{����I՝�X�G���G��w�P���V!���][f�0Y:�k|h��m��|}�O�G\��d�=c<+�� gӪ���jY�qElEK=�J26��,�wpu(�JQC��ZO�HN�G�p�X�۷�!\mj��::��ݓ��{��)2[��̺�5,�
S,�����XC�.NAQ�<�~�r��4�%>\�c;��j5&����ìd:�T�פʦ1O�Z]�����e>R�՗���MLa*l�؄}�\g�:�i��uf�Q�+�h#�j9��sf6曀9�g<���{���d��-�c3�Y�u�Z<L�֎����:����d�n28��vv ��̈́p0p�v������{q����;th%n;���P��a�L�
�PC�j���6�mN�g|p� ���#����A5�0n����Z����vO���dΧ{�"�%\�Z�8F�b�i|&�R������:�0 �~50�(o���&ZI�倃�������,�c���+�kag�<�8�����,�=�`�zUο���1��]��"Pk���O793I�`�P8k0�U�؃"[�чKl��#���!�I�,o��j�^��5G?I�D�C���Pd��9�u��{�.���۠�!s�6��Jcl�$�a}��lp�H��Z�N�F�N�Hw��
q�q
Ѻ}9
��N`i��7Ӱ��e� ��GȠj���^�K��"�)�Ku�ƘSRO�P�x�M��p�������#�����> �U>
�������&eQ�p\�e�[��ɪ��<�Y
�s�����<�~�kRL*�-vR��^�{ig�H����@���
���a��c�C��6, ~L�,�,�]*����?��
��# ����䁖������g�	K���ζ�U5��l^]�����
us0`8yg�ˍ��x�M�M���ӘV�����}��4"��犔�ZDԊ��y��z0�bl��vT��n,):�-CC��A�`���ᐙ_�:�mU���|���f���DsrVX�e�v<����K�~�����2=��ݼ�gB����>J��I��7��J[ ��<c�M�Y=0-A'�V��󫒦���V��|���1��|��4t���#�+d�@x����U8����g�n�A��ż4���\"�`�Y761n5�����xa&t�� �2@Ʈ:�,�m��4�-q��ecFsl�KwW�o���W�K3��T��(�4k��:�L�����(��ɹҬ+��|���|)��Ib
r���1j�Q�8�c��)���SXt�h�PH@'��S��B9�)�x�1/GDM��(�.A���A�$�E=��H�$���96N��	ͻW��S�&�:.MD������v?�^��ղ����Q&ɑ2f"9��[�'8�ozXzX����A���a*�����z�Ջ�W�6�<�t��N�c)>m��$z�f=to��������uȡІƁ�إ�r���Kt����:�8�?�A%̆h�����~"-�cx4�C�9���"�L��zN00P4$p�>�*
���'0f_O�Z'�i�	����g6K������78*B~Ҥ����U�����=�Ԭ�Ϥ#�>:���eY�-#�)�B��^�)��I�df���;J�6Ԏ8(3����3 H�&�v�.n?n;���t�:]��q��ԪO�0�f�i�X�J��@PŃ���P���V���ׯ)��.����)��RC��IPJ0� �7s���K+��t�Bk��,���y;�g�;&��E�1Χ���߯=�����M�L >wK?��m{ޡ{�_2ֲ����ζz�g[4��,�6U��с���R����PO�Od���N�bo@& [GXuh���I��HL�-�0��&�n��-�#.ϊ����-3��a����xi~������l�^�%������۱�B#���������R/]�]&�r�8�̹n�h����P����8��u!?��5�6O��}�u]A]o�V�$I�@�(���S�掌~�K�NG���(=��{P ����]P-ˏ#�K%���;��9��cd7���oqaE'?�WK�H�Ũ�&�B��Ql��$B6�06
���ӚC��gI��v�Ke���Q���M��) �A_��s�H�k���ak���^�$�8� �G��,:�SU��e��b1W��]��gΣmZO����9=`pT��wq� 
ҷE���4r���h?�sN$��wslҖ���i\�&��v�]\�"�h�R��l��P2I�1ѓ�0ͧ�\�y6���?}K ��S�PUe�f� E�OVy��bI��,�Չ��L�d����z��/=QG	J{Rc�"��#P��HJ�/�m�YH���F�����o>)��\F�*n��m���7P�1��9vv�C�nÓ��s��0C�"d��-��ׂL%ab��l�u������������5r�ܺ���u`/�߯��DtM>\D�'��h~�ic�%�	$8�d�^2k�O^4~��X��S>4�L�� ����f{2�o1�j�FvX7�۞���D@`���V����ڊ&�txJ������tﴴf|L!�P3һ�z������������;���6��*n�{F�;��-2^	���gO���[�+ݚWDr�Tu�B���M�Brq0�e��Χ��b��Y����X��V1�$��~�DϕP��|	u;TB�ǚd����}ۢ����N���sj�o;��A��@)F�th�'��\\���1 �6@��,h嗿Et�B�7����"*��x�V��
1��@n��ڟu
�%�o�0����g����S&���1���L��X��穔@m���րo�/{NKC���7�Я��1e����\�x��{mp m�m��WoS�������҆=����@Q.��u��@��A=�Zo�y婦M���-y�n��=����ՠ��� � �ۈ��:����Q�XLP�!��]Q[���x]
n���z���4܍�oc��m��ol�Ո�v�9ɒ��^�uu��F�kY�^�vv>��U��e�䏒m�