��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�w�tܔ��=v᫰k:����	�jQ��Fo����R��"���vE�y�DJ����C�>�>��)�J����>��4�|�j��?}ɂ�N��R���5�V1(�_�,����@e
]K�-T�����?w���{�<Wm`;GXY6��(��#�:���"3R�}X$�����Z���!� �v�֍0 �@��]�������]١��h)�'�q�I+*D��@����v�Ǽ0í�'~��@���Pf�?�������8��p"m���,�0[�ӣ,�����}�����2+�
��>._��e_VY�K�a�=��˞5�l�����\rK�#���sz�-���XO2O�rqM��F�]1rU�~��n(�X`���R�hb�
�����W��$�J�Ŭ���?~6�֌���d�����*�[�_^�j��W?���(�R�7�t(�O�a�+$�#�t�SL�����0�V�����s'�EmG#�OJ	����WqE=)�s����9}V�9�u���v*
ܧ@j&v� ��{��#��rs|��A��O��R�m�H���_��8�ۓ?l.v�2�0tLvH@p��=qT@� (�?���WCfn3��>��6�4�w�u��l�3ٿ:�.�W���A����bR�Hn�*��	�A�8��-;iM�
�E���}w�օ��}�AkH[��z�y�4Xe�U�U��R%��W�c�����Ľ��^1�(¨z�&�������3�Oy�Ѐ��b>&f*�zW�7��+1�p�7�z0q�^ɹ��3��a0�z��o���گ�U�8��Ȅ������H�a��}B����5>��A>� �Q�_3t����)f�����am^�*�Vc�C�\�YD$y7[���w�Lěc�ld���V&/e~��M���(��lz�dJ������L�R_�k'3��!�H���5�H�����}�������Bgo���()�KlA6��.��JSԃy'b���DQ�o;�}K"�I�ܣ�+�ϕM���t.���5�R�6߮�ׄ3�pN?�^��f���kJ��i����a�O)��m����=�ĕT���#H���\TcOC L���r2%:w`����P�
:��M�F�*��(�J��[A�7��ʿ���,[��Iю��d'��md{�E�xE�ۘ_����#-WJ�_�qH�\����ڷ?TV�z��5g�;���1ݟ�wXg��O�<��Ev�|������4V��'?V�>�`S���������-صE4��(ըDwqN�]�0\��6�����
��ko)_َ%\$]�FJ�c8������6��w2�0:��1�~�� B�G�F�T�wIk�<ְ���>��S#�R�H#��@�I�>5�m�ꍶۇ���;���IT
�!�Sc��O�׽��1�\���a��e��?��t]xp��W���z�0	u>�YLj>uO�ӭ��؛,D@b	P[��#�28Hݿ�Й�iPt�!ɨؘ�[�g�Ǹ��-b�ڸ�$��a7��%L�Ǆ�D K����.�kK�:�h�~msG���ne<<�Ɯo��