��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4���"WYj����i� �N�7A!�@<e�]ң�;��5DXL�%�����f�"|���\y�]d4�V���(h��_Ϣqn���RL�/� 8�OK���a�Z����IL܅T?5
�Nx0��Ϳ�7͋)]��2�� ���S-��<�&42OƱ�%�N�H�s��)}��Lo,����;��?��'[\�W_ ���������=��hm@W�)�c[~+�!?��IX͇,�ټ����C���������ۇP4��	ْ�:���%I�;�z��ؑ3���M�i�|���[m�=	[NC̩`�D,�!�>�27���FN������Z1IbR�C�4gY�#c��,�1wP�_����=v2t��˗5ʰX�v&G���|���D5��uD����Qm��ۏn���HeA�rv��ҡ�g{C�&x!o:B2�}Z��z�,a�xO	����f��x1I�����֞�)p����mB������@�k���q�;�+�Ne�w§&�42��j-��iL�x2c�]R� v;"6_x<�u��'��;.Y�)����7~�İΥ�$ŀ^�\�<�'�(�CA2���)[�u�nh"+RFa��O`��)�[̟rF��-�����r\��e����V쑋�-�냂����>�1^�<�{����;S�'��+BL��Brf�(P�h!x̖N�^H��s�"�z��ˉm���#
�����/�K~A�8����Ez�
FF�y�A��� tG5��Y5��+NT�������z",�/��"���{�}�š����ީA�*̟��ρ��[Q-���v|d�T���$�#��L+�C�2y/���4G
�x[@5N�A}k�μ)�u�]�0�N[��0%FzZ웼�&Yt� 5���F�S�.f��wI��! ��m�i���|�՞����UXWؽ|�7[��N+�p0�$ǧj���!��GJ��Nfk����J'�
��_f����!'�M;��z'��G��s�$wv	��9��Y�$�4��-�J���/�ٲ���
�e��b���%'�F�y��B� �犮�r8MY?��Fve� ��d�^{+K��4�c��bv6wj��fŘ>V܅���R
�h�Q4�^�h�?5~���!�zʵ�.HU�b����<pL����[�S�+���g�g1��V�Vr�q��g�<K�^/2��b}XgGO@}�$�Ơ��H�|ގ��}��ZGT�]���^�sX�f���⃡�e1E,����pjmܸ�_�&M8��7��UIC��ڴy���sq�sw؀���T�i�y"G�^�L��Xäs�fpc5�4��*�|��<&��Pg��(t�,��ߙ��ӥJ���X����,�]�(W�?u�������Hh��$� �^�O�|��1�]r���m��@N+�q����0j�}:�y�-�nC�� �/����Y4+�"^3v�D���� ܂zOo�w5x���KI��G�8sQ.ۆ��`]�+����_�X�#���)�i_a�q����oXk�9U�J���͜�� 6F�S�S�����%-���5C��[�;@�38�Yw��w�ùK��"��%ڤ��o�K�C �y��g���gI�sky�3镞�>��0�RR�9ґ��[�$2�
5݌�.n�	;�F#�������iUP`��E#u�q.S�C.{���0p�h��׋.����B�2uF��2š��Rv���=cɨ>��C���/ǀ�=���n2�yN�GҞ�R���Sۗ4�t�H� �Iv�5g�W��w`�܇{�@�F����Ɍ������


X� �2�����q4�C������A����Y_��d>����j1t2$��`Z�̂�*88s˔K���-�`I�g�K=�v�g���q��(J����飙7�n����w�2�v�����(47N��� COB(�D�L]�[�������~�+��=�B^?$L{:�s+��g���˗n_s�PA���o*ʠu�"���������Ko_�
�$j*2���F7ܮS(�G�j�۩|K�6	[_��c87�͆1]M�7��K��H���4�[�֎U8iY��U��wcUu5r'ı�xi;:Y�ݯ�+yڴ!�
*��g7��c|Ř��( ������@�=ĵ�L���r�	2��=T�6{�M��ΐPG/�KDS�c�Vb_�e�����e-����#֯k�D��ɟJ�?�M�ͯ_���垴v�`�� �M���Q�y���h�}���ȹ��>TRW�g��n�Dmv�Bt0�v�A������	����� ^R����!jzՊ1��i���1���v|ǳ	&=7���xE�<���
6O_F��ө�u�����X�E�Qe�"xaau��Iאm L�@q{����5�/�� ��
�e+-Ha�jO��e#��7�j�^j���h���3�e�I��〶v����R5ɢ4M'��!̠w�q�4�QJI���Xw�������E7�ps�P�Y��0}9�dH3M�FYR5XiԈE�V��#j�|j
��a`�Cr7�x�،�T��%F����@Z�f�������$��~�O��ֵ}Tʹ�,�9�g:jk��q�6rR���$ճDd$��ޛ�%I@� �h#�Kht��BF�����wU=�y�#��I�m6��X��u~i>�ª's���=�i	Ԧ�8���v�D B�	*d����=O�n�\��K:�/f�JDu�|�mmE�|I�D1a��TzM�<��o�q뺊�<zL�x��e�}��5��~�#�5_X����]�\��,s6�JP}���VQO�8��X~X#�V�Ƶ�y�E�(%��&�'?�,���aG����o�]�A|�]v����Ԙ����U�yt�23�~�aɜӜ��mzѡ����|j}o����i�4�ǵ�Y'�:��e��a>�l�h�_���`�7���C��Pd�<��a���f7��T�=��q��o���N歁���a([�>i�3�R�� ���{]
v�5& >�m���+��.X�v�o�J+�IK:
3BF���|��a�5����T���T�B��N��]����+4Ζq�m��8�9���v��ڶ�O���n�h�^��Cd������23�*_�Cx��J����U��Ip{b�zk�Ɛv��8S<����3��9�f	�je���e��RS<������F��y�?��AQ/B��t
�]'���Y�T�qz���Uߺ�@�u�\_�x2p��{�j��U|�H���I%{dAW�����#�B�/������[lscI3���^i��@��ƽ�@�-v�(
U�,���Ɇ���Q���[����z��c����-����bb�(��+#�=�[.�'�8vc����GA/��w
u{��(��sy�F��YB(��O@&)��y켦�2�Km�~{*=#�ݬN:��Մ.�t�h�ɷ�<I�X&�\U&���*))f�|��Nt�A���c{��Rr3�V�\ �P�H����ViЙ5^)�No��q=��m]�ۇ�f�`��A�>Tb��m�c��禸'=��?����x.�.��JC��.0"���ڱ��lf����r����dc)�Rb�g_4�]�$>hb�46\6��������6q	�^�ͬ��P�Z���T���RBq��'��䂎�;ټ��et�PȰ���Ud��xw���F'�O���u&%����@���t?W�E��o�k/Э��+�"�+�LJ���*6��w�1D��Ӵ#��Ӫ�11��sN�Hkґ��<#�r�{]��YF�
�`��
�\�{��س7�H�k������ �������/ �,WZ���/!;�M���c#ۑ��eh(35Q�eݲ�ruo"PS��Q�W�}�� ���c���L#�X��5����UM��uh�,
����W�;8���O� ���ֿI��� ����[�������u���rޫG��q�SR(ܩ#]���hx����y����7�Rm����ŔhI���t8���h�p�L�]������#u�mj���t��@�.6��:O��~P(�g�|�o�)ڜ��`r�_��(�8=�'7�G�1�Mw.�f����va�Z*hMi�o