��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�7ټm�lQ�חY���f����ɟ���ZXg��;<{�&N����~F�x�	�4��Db{K�9�n��i`7_8�@�S��T*e�4].��SP��ܐ�A�FH%��m��8��ucQ(ezc-�.�����@��
��^d���v��dꑠx���o�A(wL�q������n�"��H�Vu�PLЙ���Ձ��'���i/����O"!X<M6;N.�%��a�X� ����'պR����Ԓ^�>��>���� ��ş��I�C��=Q�/�|T?��#M�i(�z �D����lH���J����h$n���A�qI�Y�JkB�˲݊�����>�zQ!p�&�x�]��"����/s=�ǔ[�9�;�7�P�����5�I��8�� `y�gf��qX�1�w�f D)�%~W_�)J��'��i-Q�����:�<��"ԱoFT8�3QOE����a�%�;;{P��O)�i����A$.�g&6���(2��3GWtr�ZW�@B!�%RE^X��eH�<f�MW3㵽��������fK��"�4�k/Q�l.|�-�	�5&�`��S(�CԨdz�3����+j�_��ƕtj�߲�U�G-)%�'�k*T�=&���4o��%�ԑ��|K�Pt��F��_�KW��R��ObP��J��_Oܰ|��
˽���i%i��!�թ�tYv8��BuN�cS�M��z)�3 �u�y�i���iqM�-�|�V�f&"�t��Nh���N��?: e��+�, ��L��bdE��0I ��27�"� .q���/�<|m�+Ίː㹻Bֳ��a��جbz���ĉw^���W$��	�oU��^/3�=���c�K���`+B<�ZQYA���`��kO>�(#��m���!���L_�""dt�SC�t���cK�j0�E^�Kh��ѧ��tY<l_�	�Ǿ��&ǖ��(��/��i�qvo�G[+W�?����0D��%�
�o���7�N&&�#鮊&��w�]���� �SD��n�/���=�}���!�O0�����zR�4*b�F�ݮ���Ĕc�5�_v��k����H���d�4�SY�s	�ܵ��'��8#���^ɓ�?���K�k�80�
5k��i<_���S�����s�8�h��?���SC+����cl#FQt����b4v�F�(C0+l)�@�# �S���嬾f�X߅�w5��c��/N���O��
����E��8t	i[�5�~P�oE��wLjn�i8x$n~���vϙ;;�ƭc�V��T�5f�5�����* �g���k�K{b ��\��0ƙ1��|4������c�C*��˾��������*����o�ٶ����)�%z�-uz_��x�@4k;��j:?�۪0��%{u��p���KΪ�r��{p���I�42&�q�JخC���2���hH����*Ĭ(yb���-����'��JL���ft������RY��!���<-��&lT��1G�H`Ce�߮TώE���Z�D�M ��<5d˱L���IS�N}�; ��b��4T��H�h�݌������ ܭ-M���t
�{��z`9#zZ��w��.D:�S〺�w����(8�-T�'$�ۉ��h |	�%���;֮Mw�B������ŽKh�D�#���K�t����8����Vd�`r�+�3Ӝ�ԅ��c�
-rMF\f��/'�L�hA�I��İ���h�����N��O�(�*C�u淉T�}�9��l�"�����H���/5v�:ɍ�gx!d���?
�j�����6=�h� Ü���"����t�=�L��h�Ɠ��n�1KK����e8�n󉛶��_�G�MN"�:��=�(m���� �����H�⪫��NR�� ��T�1�H4a�|�Ӯ�;�{@S�4Bi�Zޔ	d��k�X���id�^z��`�����[8Lv�?"�IhU�y�����0�J"ߐ�� ��Z�4��.�C~�W��m��nN���K�ߋ�⠨�̾퇇KJѓ/�|܏e�B�_L�n���O�PNM���2$�܉ftNK�@����s���<�cQ��R��p)k�h�E�q�f��۵�Uy>(���Q_Έ�P�K2��z�)�Y�q/uk
�Ī�r�gW�1�Wh`��~.�PB���m|��Cz8N��F�i��	{^ǃ|��G�gl���f�LN���9@�im�L״o�OGw9��J��e�L���W7�m�G蹜i���L�GR�}���1J���R�G�OD��]���L� Z��y1��b[d{����K˿]�Tⵕ�y���r�I�ݓW<��aNA���K����Jk��V6#gq|�G�?�9U/�N�.c��J��HK�
� �v��� KZ��VF��|��l��K�U�|�b(T�W�	$�@s�R1V��?-k�=U�)���q����F<��"�zLp�I�5�2�5��U�$��u������m7P1�PL� �l���W��I��!���ԯ˜�NU6�1q`��3]&�?V���	"���"��w��T��`���3�#��w�Iq�v���3A�Պ��{��w+���1{Sn�2�؍�͋�\�^��d�����x%|����Ͻ�R�Uo�	LĐ�FU&+��n]��,��]�R���J�}|���unhF
��Hsth����w�:~_L#fP�*+�o_�9Ь�Jq��/��Xmdm�����[	��'cCmE�;*�+���k�A�RT5=��.r��k�)�]k�{LH�I��xLzؙ$�۱�_M�3��xą�▝I��s��w�h��=�W}��Y������������(�J��G8��||�F��[�XF�`aFJQ)(zʳ�| �