��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P �&���^H��L�.�Ia��@L`2�`�̗�[G�yu�S���,E?_�B�l�ch�o������֝|�v-K��������
�^'-<�La��U#S�9v{�Y�.��ٍi�	��=@$Y�6W�:�m����@}&�����x^��Q�	�� ڥ�St���/=������~E�����;�NjI�릸�n�R���:g�CSeѻ���l���bt��d�(�&�ه�DZ���G���qٺS�{o�M�dE��f����:o.�B�2�f�_�u�S��2�ۋQE��
�C6>�(������=����=�ys^�e�[��"�p)��Pb~(�k;�$S�U�c����<f���A�I!Y^VI�V�����Xn�!��DBi�q�<�6\���e��?�_17LB�q=���~c���"���;!��!ُ��V���`��W�@�ڦ'H蜧Qݩ��<���ǜV@~i�ro୰�.{��pk2�A3ѡ���X�7�ҟ7����dPY��u1�J�`�4)��8]�ՎbPeG	C������s����W/4l�bn���?� ���Hf��c��M?�@�c:˱��.(�	{_�x½!Rq]��Ԃn0A��*%p�q��BrAe-4�sx<�{���f.cs�#T�Q�t���Q<"$�㑯u���*�Ș:����~_��1������W��
:0���<�����ԝ٥���w#IAX�g8�i��~S��N�};�P.>��V�+�"逸�a��Q��oӾ�[ ߘ0�*��n��+�T� R<�qZG��� ����o��(Q�.�Cm������@��Ut�ڋ�o@��8��Vp����;)�X�6�~�9�Q�|7fj��D�� h��;�����g�:ǋ�I>p��N����	��2+&m��uX�و��كM�*���y��A��NT���j�\t���oQr�y��U�j��x^�<� ��ؚɶ�F�%Y}�����<�)�?���΢�D/���ơ�")jii?4I��m�>6v٤}TxIзP�h���u�=<Kw�t�'$xL�[4��&X2ʘqγWS�T�zBD0Y� �ӑ��OH�D�Y��.��p��6�
�YKcV����@+�U�˙B�6�N�Rw�����T�ǈ�p����E�����5�ާ�4qg#R�E��Y�흚I`P�, �r����:��g��2Q����콈flĿ�t
蟋HyF��,����������S06u�cMT+jy��A1ɞK��b�8��s�~���d��Cƌ���k��DA+d�@�k($��0T�n
��a���(���';�G�}��Z0sP�^��<�����I;oW$�v�����l_�����8ڶCJ��þ,���t���v����gb���ѓU8����Er�z�a�@��[h3�qӳ&������[XN����Ox�k�:i�#�Y���떯�LS��~%�[�	u~��3��F޲@�>��a��%?��̎&��$�b^�b��0���J	���Q`��j; e�]��<�Z�ދ�#k{P�@�t.|߇dh/��`�mǰ� ͸�>	�da�4?�e��PO
jY찼X������6���/�uF�
f������'���=t!~��Lm�E�=�ͨM���&�T	^7�<��R�)1E�{)�p��x�,�;�����<O8��x�n��"��CȌF�
t�|�"%hR�R��s̬�AD�>�gu���<X �K�ی�Y���I�3zdb�6$a�� "1�?�Д7f=�mq��P��_;9���$wʝ���l�v��h6l�T�z��6:�(�H���JXUX�"N��R�⫼8)Mt߸ԾuoOA���yM��ڢn}\��M-�{��:(�yZ�w�M##߭�l�0Y�)�,2�<�U,��Ĭ��-�N�Gy�3v�]�?���r6hA��ѻ����N����5Lf��?�T�"KeX�!�UX��˨�Tl��n�ȶz��OA���3�"㯿|���b>�89TҿƉf�"uJ�L������5��G|6c�Ei�C2���U\DquɄ5R�\��K�E�E2K��AX<(��KGqf"�
�8�y>�:{��!"�����d��::��ֻ�"a��u�{'�W# 5Щ���%߫j��]w���*��)�����x���9A��і�s���k��{�eS['�:�s�x
 o���f�C�
���>g�T�(�A��:���ܟ����_��.	��T��?X�E��a������D�<A�cŔ�Sqo$�-!ص�����q_��r�q2]`)�$�����(�ϥ�Y������Hڦޥ�U�H<��:�R% �?��6�����Q�P;�êU���AH����|��ehh��\Pn���2�9!���Wt�.�3SׅW���W��9̛b��Ys�l��5�{���4�g2(��e���3CNMy
x�x��q5�vK���jPh� ��H�#"���B��pP
��9w�V�����-�:���<����b�hO:���_P��hU.������GPB`���O��Ë���|�Y$��=���&��k
ey\$���F h�bX�x���4���r1���vv��� ^H�y�0}�6Ѵ?>��=k~}�lc���l
�:�DAa���M�o�['��c�&SZl���3�xz���k����nD�� d&�F���5[��R�.9&�H��G�VS��k.ؒ����4:)o�٨����B�huR�f- Rt�\��u�l�m��
�Ld�ւ$o�e�z����;l�0TV��/�.J{�u��߉P��(I�WOVӐ��*+Ѳ�/Ϩ�9�j!�e���Z�i��c$y$4c<9�_^�r6�F�r������
���w�O�ſ0`٢�z5;�=����-�޿w�
���t��Ӹ@0��U������x��ߥ��5Ag����UC��I�Q��{�E�\̳�#�vW x�Y(��q����J� g������ӢO�\&�d��c������sY������ G;�*��:Ê�����cnL���&��3�+��L[_��/;LpA�u%�	`����W#�Ug=���yf��IA�0��Wx���[��e��L`K�+���&����m�a��UW�Hg|~,C7��5#�mJ!q07��d���(�H]K.��Z�u�>Ew��p�t�l�L�R��X��Ǥ���@��g ՚�WxI�b�?k{O���������pU�7�T՞�O��U�a"�Ob�GWoh���t�r��_�:+aZ��v0z��8��A��˥��!����dk�g�č��_����}�Z/��H5}�āTF���W��0 }G��c܎3��t-T�[��.���dj��K��g*�r�R;�|G V��w� ��t�H��t1l� A�:@*��2��Q�.H�
�߃Ef� �i?����+�.ݭa*��\'9ݩ��c��$��d-�k�/Z�~U*(r����{��2����� �"b�>���?�#=�vy�����D�b�L֖����3�w�&���
{I��JѥN�F�� #��n��U��SA&�Sk�:���bж����}ʲ�sG�(��%�C�� �s��t�;Hf����=�`��:I�b���5ЮK�r��sN��u�-X?D��q0��J��߄
S��o�Y�>4`R��ͪK�Gu��/���l���яv��g]�������0���/�҅K��n����+ܞ@��)!v��@�������O�*��#b��q���kR�ek�r�o�
kc��^VVo*'��k�;r�Z�[1���-~��!AaE>1"I>��Z��Aʥ��s׏�-p�F��B$�"��V�����~}v�_���ЬL�H��_��BY�[��\b?�Βh`������iK��9�+�ܾ_� 攊�P[�o}� ��m:�(�eDN�l�BBg.��U\�����d�(�o^��@�"�ۢx��[Q�|�MYɤ�NcZ��&܉ږ,/�
�JI�K�VV������o;�^�{�!����&���yؑظ��ڙ�@��^f�`��Lxp^�	*-TB�}:fH�ҍ�Y��|{Jmֶ>���ؓ��ɖ��c�M]�ȑëʕ)� �۫� �z�_!Yr��-R�0'v����7&��H	D�i�O:j� u��r�qB{&�F�\��m'�h��"���,��V�4f��C���m� b�bJ��WRa���������dyC�2d��V�#�X0��d#<�x��M6r\��\\xA{��zIݦ�Qrq$7.|�L��,�p0�Vdp@�"jnj��<c�Ȑ�K-�"}Աrc��([�zFN`d[��p�����	ezk�-��G��ϯYR���*P16�a6��W�Ů��C�锱P��^�$�J��*ۛN_��Rj�$�Q�|�����oO�x��v�$b���_o�Q��R	�v/�'�L��$�Q7������灣'A؆h�f��i���>]���<�4��I��bEcW2ǳ��@FI��o���v�bü�P#佅��[[D�vD˖�P�� ֬g�Ý�C�g����/��j��5�̴vG���Rg�mҐG{�kq�n*��8��~2u�V�� m^��Y���G�W�jpo��b�)���5x?�M�a1��OD���]��Z��+1؅��(�Zqڴք�����#����	�q��ʿU�D:��8=�JJ04�!8���j�ߍKxXm�I�=�/�����Е�V����s�+�`�D������):��~�
�1u�Ma��Qu
�2�Ad�� �{����Ȏq,�}Ly���/����`&@�s��B5�R�Y,:�i��6*pμ8LT��R.xi��y�d0��yT=�������`�Fcj7��C���8��� �y��ǭ��/`�v�v����s�>�j���q�9ｧ �+�����*ft�C�B��4Y������b�,����oҫhŊ�]'Uq>�9$��Ǽq?�d������S淺0Hĭ/�N�*z��Cd��
��М��{DT�֤�W�^�3���3�6���7Ι��]�H��խ�48t��7��Ь\�⭺{�]J�����0���I�|**�8Q3;1�M=2��RK��� (�tc�P���i�� ʑ���Z��cX��̕�	k�;�����pMn��$A��-�,�Oԟ}�������:߱��E]t��GVn�8e}͝�����=��	3,�چ��j��2ǀ��TO��#z�.+ww �_�m�����X��ڞ+Z���iL�-{�-@�2v�*߱kj�[>��=�u�IE��n5��8���8�9[ƴҋ�k��wFy0e���rV���t�𠳔Ĭ�^t
&5�y��?�*#"f7,6��G.���2ܣa�[_�j�� ��71���4�Q^��gOkI*��Nv/�� -. p����9���K!�W?Er�x��s(W���n��(�D��/�%֨R��}0��A~u(� �2�B��ɬ@�h��d�*���;�*�	���{�p�J�6�xg�8�5�mDwu�{q��+���k{t��ò+P��8�L�9m��y���8 ��61���Ę`�M�����BC<�N�%�Lsyk��[�:�~���TK���W�;�yq/L��I*��9q�-i���>>̊.��FH�N���W���Z��]�V_�v�n2��*l"��v�G��\q"�.?G��G���'Z����]�N 5�_%���b�v��%\�J�ԚC��s��'�pF��!�iB�2���[ܶp݇^��y�Z_x/i'~���tY�oB�g� 2�)�cK���(�h)B�4��Uy6R���O$��+~�6"@�q\�����N���b1����5HX���H��@� 5�����y�jh�ف	*h�j�H��S�Q�k����ɧLT�}�_��ɨaH�� �ω�X������p�� }�٨�Y�y���w E�u�~��1%/�M��%'mOŬɀ<<����C�.���<�=��u��Ľy�윢3�e��xH�J�~�x��V�FS�Y�Rs_��n�ux��S"�3�i�1�Ħrb��qn�RR#�"Z�_���(o���O�r��!qZH`7��;���~���Q�L �]V��|��G�QA9'lː�
��]��	d�)��`��r>��.�,�at_Bv�" �r�h�8&�r�gڧ]��=~��a�ۏVڡ��<�ւ�762�%;g�B�!\��:��v��`��q�D<�	1�C�i�"���<+�s6qVR)N���4�zf��]��A�ٞ�cȤo�o��;��-�l�ɵ �ԗ����x�!R��N