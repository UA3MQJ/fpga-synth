��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>���q�;�;�g�?�_�q�-�m��5ʞ�œT����
��cFZ��R:�'��o�xE[�I�N���B0ˀ�2|:{4�C[�p6~��n�?�Ϳ����^:٘�!,�i�dF��<<���0������� �Z�=+C�r�.3]rw^sJ��J1��`g��N�X_Ac�N���W�o\L�(&�!W��.5N5�(D�Nj�D��M�'/@l:F��a9D��B�g�����op\3�<)p�e�Mm?@��¢�aբL�@e�A�,W���J6%�@F�~�bN5k���kh.�t �$���ܔX�@M󋶮�(�
Y��޶@�c$_9�e�Iߜ�ui���K��U8��6���V�ve�Z?7��L�¤�O��Tm���UX�5f�@i�?v�B��>g[�V�Ꮘ�x��!K��͙'ۧmb�]ӧ��
��#�|����m�h���%��'x~ �s �̇��~��Q��
Z:�O��+3�ٷ@2�!�$}��{����td��0?W7��9y� ��;��m�rЍc�ݴ����;��������Ts�^6���]��s�_[P�?�X�k*��b$Q�@�Z�� %v�J����1>���C� \O�O���^�f��%���Bw��>�V_ً��9��P|B����/St��d9�z�����*�s��ߎB�O�^�!W�� �F��!����5��3�*t[��܆��kRgSdfAi�_z�Q���N���Gp%�D+�`����k^~��X'C@@B��̟�ȋ�J}�F[E�-�����.Z�Q���Gx���0�q��|�{���
�d��sj��3T�����|��&���-1�f3կ64Ů�X�L\@`&O��Įk8�T����u���|��-.r�"������]��߷�ӿ3���!��k��Y����Z1��W`��"*yR;�A���k92;A� ���/�8�I��S]r�ޜ�@�=��A�ő#T���R#��a9-�K�ө�_S�.ɚ�X�p�LO�=,9S��W�0�s0d�p@.���k=�*�Ax��D��*J���E��w=e+$>-�&ۑ�	���	��]�e���n�������װ��-H)�#UM�k����?*�D䪫-�z �V�{�iK��(�J�l�G\����N�A�HT��f��S7�{�,:8��!Ik;��}�D��0�NK(S6`��~'�PGt���pp��YD$�P䂥EtKH}Ɗ���_���jٌ[�.����ͷ�d�^H@��R���iB�7HTw�`���y�Tvq�X���n�%���"�c�?ؕ��4mEo�Kc��mf�sc��Ok��H�2To�)zȥ��؀��I��gN"|{f�d����{��h��.��g�@_���/n��B�/fby��@�c�{����>P��a�4 �1�Vn
e�a���1AO@�����(�9��B&	 ���_G��(�B.�{�����W���u�T���O�HP�޻�`Z�!X���/���o�a1�rϖ9��\��2��L|M������D�(��z5T¯��[W�k�� ���FE�>���ҩ:��b����4�<����?<ܭΪ��5�H(T���;���z!e�y�����ꄋ���`$��pĔ���qp�2/v����1F��?��|��q�Ի7�$���=Xo_#n��4�_��
W2-=�K��Oټ,�vM�WPJU����*�"�a�7�kU�H��zHU{n����9I�i�n`Q��ǈ�+�k��ge��\���}M� �=[U�x&��;K�FZ���?%�͆�^�Ǿ��}eo�l�����QI!û�,~�"�b箖��6xv�E�6��`r��3C��K\�vf�w����1��R��'���1���W��$)b��wf*|jG< �#Qj��di������qeҾrQ������\�54}�E�VQ�{"� ����y�k�F0'6����k�A�U�R�0~8�������
��	�lͯ0������6fQ�D;���eixW�ûz�a���Uŧ���8J�,qZ%��Gkn�>ѓ�/���%�Af V[b�T�����7���/
����6u������l�Z�w�ӤJ��ak���v�&�p�iC��z���	L�y��Fd��`�RO�� NRQ�t�����R�Qh%���E9*�p�Q�u�|�Co�^^��l�gQ�I�h@�p��+�P�c���EM� 
� ���7Kܟa�Zh�G�nt�Hé�t��h����<����4����ln(�"��3&�&�i�L��O5�U�Up����6&�*y�8���ݓ�/Mwu��n�6d�[+�+�k_��x�8�x( �~�E��Bgg!�"��E��+�w t��'�@�5F�*��f��W��vQWǄ���i����ݚ��#WZ*iT j	����^����v0H�R�3�Ў~�� |���V������؜,���zz�.8�~��)��+�1�	j��ԣ�S�j�eb�vl3ׅ7و�j9�Щ�p)vY�GR���g��_�Q[�L��7x_��3�i��A����Sw���;�HCՀ�|���ٰ�jt>Y
/=�Pҵ�zඹKw��y�×�ʹMs�4/�)2J��m�z��!]gT�r�-�D�,{��Ɉ����r�
�>
k�Z��~��]�qܘ��g_��no�B�p?��{�0���aN;PZ6����:=�-��6~-�rwe8�_}R�������W�&������$P�k	�e�A��ù�P�s��v��N�W.5MW3�*pe��e7�&���,'}Mx.��`�.ω�,�s�WQ��W��3���u�gz�EA-�[BǍ���cњj�{E진cz���_l��AO�|.�b��Mx*s'�)kS�Q|pR<�hA�8�vdp}�z׊�I;���Xb����=�8T^{�^��,Ӯ֏�e�*5��kuc�Q�*!bE?ES�Q��1էU�S+���vK��{�/6���zg���܂q�=�K��W��D��-��Z.��ႍP>CN�h�;WU�\�q+a#�(���* XzT>��h��jbh�J�POz�s�`y�c���g0�>N�;ӯ�M[X�Q�۾�Я�3�!�W�B��w��f�m���N��|��R��.�l��-L�cĬ�9�5{�z(��6������C�,���_�2*�w�*�o��z��-�1�@��C#�_	-m��{���P�i����pD�WW^}��x*��.=Qz�4%��KOI.�h���]���3׎�x�v#�s�vf�B��&gu��xߠp+[tp�N�B���z�O�s}��s�t��R��`?}��H��aH�x����(��.Hf8N �e)���lg�?����-�;A�[���ҾV�a�.�5!�'n�%�����Veo/����0`E܂�C���Aa�(/s�ß-�5�,��P�3�F�>xw�����V7J'���g�tH�H�f�&Rwԗ�DA���k#w�m�[�hc���[��u�"�i�M����wP���:A�07ɓB�L��l)��w;*��*nC��l$�1M��j�v�e�YK��2���n���bɃaH�h�ձ�2�����O<��^�Yo&�B0��S�rJ���*�G6L"�ܓ#y3-ѕSL�M�]���p6[�P��sw���g�|P7kf�܁�1W���Y�X�G�k�j�"u�RMڮ�9!��&m�C�x��yE".wR�nQ�g������N���ޥdx��	�����t�9a�7"�~�$AQ(�V�"�Q!%����k���Rp�v� -IgŨ|�}[���/��~(�Ϙ nn�:�����+���B뼩S}پ:l�My��;Vx����HWI�a�Z���2"���5k��C�-o�2 ������p{u��z�9�Ȩ�Z
��W_��j��0��H?�e�����MD��G����$\Y]YflOH�͞.�*f�p/n�/��{�m[o�f�|�bk$�������ަ�|���!���c����2�����A ���
	U��Þ ��2\��}?��?Ϊ���/S��Q���C&ـ�V)@���^cd�-�}���$K>�^Y�z@$:��V6btҳܞ��+g�r�������99���~��w6E��>�hC6��܊�6$���:�4ԁ�:J%k"M���sb,O,k�n^���)
l���1��~~0�k�;�.�]��{ ʝ�4r��hxM���"!�z��&Y�鞪���y$����'���~Nr
׼��:��<�l�ҝ�T E�Xp���:P��2��e�5�/9�.ĆTM��藼�U��a��$\GR���@��G���v�Q��n�(-�����i�c��g���������0�e�+���Q��|+w���1�&��=�u���A���d�֬��@L&�wH"�%�ϛ�g�\�}z9��I"��4,�߱_�mQ�{�7�S�ۻ�d�d �N��@�HK4h	Őe�;�8��e
hi�u/�oҵ��+��`���׆!���KDK�LB�;��k���c�Ue�SN�U��'6�ۑ=�0��{0����?�aTje��љ�tz�a)��tL���?�>���{��␨=gm�]���Nɬ��%�����çyD�W��I�ѥ�1Vꂰ�����1�&�jXEVG�,���36TNv5b~6����X- ��"��"�|��}�1�,H�Hv�r�!��:�GT����ja/�٠�����Di�H]����LGp�=	<�3OP����ov�p�O����T�*�����B��]I��&�C��`��Z��ږ��f�����S7�\��;�<e��*��E���;��KRc����^��Q���}��U��IR���`FzY^���z��B��:y�9���<}-޴k�,�V���2 �������[U��k��_F�[��Z��"�p���I������,�R������^����_���]N��I���K� ���o
e�`�P��t|��*�s�=�Y��cxn �~ ��tu
p�\J�����$�(=��뚮RM�3X�:�G��~��)5�h�m���'r�#��H�#�36�Es�V��)� ���!�&�+o���a��6��󾖊����>��!gM�Q�v#fDX-F4�.?	s���.�,��gPظ�
�5��ÎNO||(�uf��i��[��J��p�g��ِ��u�� O�+�ؽ���X�Z]h��3��wl�(�I^�~�ݨ��|�q 5�H5��S4�����X2�ZQ�O�>���0E+_K�"yN3� ���ґ7����_�p̈́��r�+=w���#w��R�t��ߟ���p������a��������(z����������;�3�1��"gr�!��\P�Q
㪠��"�fbd*P�������q*f��Y%^��G��|$:Y����ꇂ����_z�H³ �׎�@�G]�P!�65��hb�����uq%�M^���K��$_D�7�˭�2��/����1�7f�����euATZza���s���Q��T�dO�������%��F:f:��5I�Z� )��6^�^�h�^��8�D,rX�LA`�H�2����ñ/%�C��2S�o�,b���|^.�cn͎f%`|�����a>����b�e/̡7+d�g��:��/�P!���D���d]����d#p���� 0��L�Z�x\tO��������Ҟˀ����K5h�f*B)x�g�fv���]���:_#D�Vt��Ⱦ �g?b��̄�*��?Ct�#�\�ż�$>�ʿ�F�r%��3av���'�Iź�Ѯ%ݔY7Yʣ�F5bF��1�Q�/�9%8T�َjpj��;�1��5�2���HOjX�[Vq��C�0/4�{�=q{ �7/����N�����n��`�S�T焳KL��6���(�O���x��W�i\�����P|{P�N-�i�+8鿞*
%��5�w�:�g�N����z��)����.M�7)��V��픇8\C��ğ�'�,m�%_�*�l:^]vk�{#C>�f��=D-"6����[(�:m298��y$jK���6�-���N�j"���"Mӂ�#�迫�,���
�
��*<ߺM��{�� �C-
��<#G�kW��j탆P̽. �~n,�a5�iP5u�c��lG�5!�1��m4�C��aءN���*3��׊�"`���kJ 7B&��R��<z*<���#�G �Ǆ[���d��������{�E�s�5��Y��d��z�h�zձ�Qt���ZG)�A���>eQ:�t�Ǆ`��4#�~ɭ��thJ��p���K�
s���N#q K
&q�p������MAq��Ʀu�.��Ϝ�i����PC\F!��V@�#����gI�J�jhfR��?I��nQ�䐠�U��k��`�k�����ɱ�dg	;f�c�t�Ia�K���k��F���N���)��^�_٣�P]߰����>��Ut#�%<Q9g���YO�,8�9�Y���:�3j𐕋�lq9�g���j�І�k�K�9XB}؏;��m��N{r��(u�^�]���j�S�!TWvD���G>690%�T3ϗ6��p�glb�en?4y��-^�����D%�9jVlN*h��=�I��*W����k)_**���nyd����D��.a[P�s������Q� �g���q���+h���Ա��.Z��3�w&5"�Uj/1��4�|buf��U�a5��t����7�O�A�K˧G� F����n����DN�|Ⱦ���Aw��'����:�	���ߧ*�a�Vq�� [�~< ��[�oW��_���x~�~y�/�� ����8�xC �s���\/.k+%&����s	�����.g��#�8�F:�gYܼ
��i�
�𤘠��<lJ�28�c�ѴE�.��q$�e�ѸY��Cmm���7l_RUZ�/��؞`7!��c2B����o>��9;�Dv{�����ӟǭJg�r�-��,�-����2�	2~�;�/]{�у]Z������H}q���s?��m�u�DSȿ��D�\�h��h򻵾pw���	�i͙��!db�(�ǹ2͎���H�S��ӌ��1}��9������D�{(����$m�5G�=i�!X�?�I2x6�4]����x!:�`T(ͤ*��w�69����>\'��91��Dy�4�ٽj��Xf��qQ\F�&���:���ʴu��O������8<|�l�lɌ�I�X{7��n����Q��~�06��������)I��Z�	x�nk*g"�w�>��f�į���{�YZ�ښ<XQ��P��Z�aK*�3��4F���C~�A��{G����
��U�5��`��A�冑GR�H�(,%�%����#��w���&	�<\.]����ķ@���sPPE̖�ӁNi��tIxzr|��JB�{#,�~>ڞ�2�s�Q�Ԡu��i%IS�`N�1��tD��*��l��;ʦ2����r��60,�{-�G�\��}v�S��*���:�;O��UKݭ��$�$���/����y~����7�+�4=�fy%��x��]�F4V.���eZ�{����x�CY2��Ϊ}�[4������%����u�4Z�@�T��:�D�rJϢe2E��>\9�j]�a�3hF-+-����뻿�V�X�玧j`�ѳ�x�vˡM1�*�]3�XWjn�Dge�.�3��fM�J>ػNĕ��S$>����-8`d6����S��x�M��4 Fk��wwJ�d��I�q[���;��IP~q�7��Ơ�/i��חZ�`WI��G�y֗*�-LKr���HL�(赆�)M���������.��9T�A����`v�A�\z��%�&X)�%���/�^����[����xB�̂G)��=�k?=�1��PZWz�����Q=&�Ã��zs��hZ�KRkNI��OP0��G��ȃ̴�sb�����|3�y����y4���]��I���<l~UG`s,e�:,.��k��n/D6��*�r��k��H�L�v�oo�m��)5�l�&RgP.z60��OV �V�'q��#�׉��3.;7�7�K�쓶���'M*4�9 t0,C5|���G^�����ý,�7�e�<�a��k��	x�0��a� YW�)�)��#�g]F�[!���"CWq��.|�v]�F=h�F�h�{v؍h�#r�Ғ���95/��Y�+"�W��r�6ו}k��7�������2��O�N����`G?��Id��P<E���(�C���ظ��f+gڧS�p�x��&.��j.�osy�%>4����e,8CSz��U�/U�q<��'3C�t�˅F������;؁ jՕ����Q9�ǿ�j"��ǁA������kރD�(݆tp�k1J;���x�O������8�|��Ov O1��"��ع֬��
.�ԝr��To���
��v����ͯ��P;�����Q�	(�"���9��ϖ�]�%Y���2�)��4�K�=L䮝V�a��(�)������� Ӱ����E���0N'��ӽ-�$ۛ�3G����4�	0\21r]�2-JAZ7�g_¢����$�6�O�T��b>�t�Z�]j���v��i��O"[��aE%���������å��qK�d���RT�L-v��u�m&��X�kU[���(f�a-�8�t�����_x4 ȯ�П�&r6�j���-"s+�t{�X�L�.>A���#@ԘrŜ��K���T���ح���X=�G�����H���Ze#R�l� ��<a4c���O���qc��}��h����7Lr2��ߘ�$�u���}�,��ͯf���T��ibt���՘^_�أk(�o��ѣ����TKgҬ�hb�6��W��:�~}��{�����&�6}����mfr5�u�
����j���N��;^ �@끼W�a�����f_=#��}ALj���/P� �t���$���:�|.�]���p4��@�4�� LSC,� a��_�P�Zg54�qH"�
L���h)��+�EZ2�1�=�����
%|��
�ΏKMm��t�"�����M�K�<�y�`�]Q��\ʈ�/���c�f$S�����	�'��	���q��TL(DD�����J -��=׊�
��ۈ���h��>�R���nV��/�-AX�!�W��iy��D�_���ɻ��{w��u���)����$�Ђ4�V!��k��!�8����dGh$�7�E���Ǎ���V�˟��|��H��5��������3��6gǡ84��[�q�
���Ȫy�	r8 �����	:�,���X/k�л��I�P�߂�ӈ�	 Z�q䑽�:�8�?x1�Z0N}�k,��� ����h�a�Q�|,eK����fF�>� ���-���0�3��	y� =ţg�&ն�it(0�5:�m����7v���{��q��>�'IP����g�,dA�����s��{~�e�>�<�&��#�;�����~��y��I'sw�:��f7C�
��"��=����ve��Q�Xhe6��9�qMew�.�s4jbʂF�5�i�`q�d���  ��p������Ң�|��� 0Bp��&[���A(Ǒ�(�4S�6-}aGB�*�|�3X�qw6pj��m�}P'S �t��v�o}����T�ű���u��&p@9�@�fL�E����UJ ��G`*��<� �������Mš����X��[��9r�@#֥W!
G�C�wD�v�4������w:�2�"$���_�r�2ndgg�4ɳ�{�#5����8@��4�,��D� n��'���=����r��G%d�~k�	����X�"��m#/-�)���ܲE�(��[s��7
iy�h�q�������F�T��� �[2�̙�Pz��O�ߧ��OT8۱��!�-�(����}�\�^9��Ȩ��oe�79Rܙ��ǀ����)"����:��޷&��׎Li!<3ٚ(g���%z8��.L*On�M$�t����;���\��HǄ-X]b�֯�/}<[{{W���ע��w�4q9��7����(M��{��������%��|�6�K#M,���a%�C��C
��Z9*91Ж���(��|�P!��&�M��� F�w`�,��E�!v�8H�����s�M|fj���|�D3�S��ū�V���u�7Y�m�z�U-�ڪm�X�w���)gFi�C�&o3� q6�&录�ߚuq��,��W����<d鋲��� ^݋�0�����M�m��C�g�%�RWX���J��P��8�6
z^I��Z����=ybc4i�/�����#h������風�_�u�1l��Se��3�<��LMΆRL�װ�7�+���4B,j4�S���Ca�r�gENQP?x�)��5�	�e��7j�����G���<�ꂃ�ƴ�Q���`��I���͹�)����{���`�x >���i��s����Χ���t;���o�Q���az1�T"�Xgo�_��ȕH%X@����yT�Dv�/cZ�b��P�.�h:��i<o��1i�����m"���.Q�;"�	��e?7����4F�gv/�ԁ�i���7V�Jj�O�R����x�RO�aS&ΰ����g1�N4dU;�p %J�A��5� �x8�)%1�Uz���W�+� ӟj���qFn��ί�R�8�xD�\��=��y�1�_u�a-�d	�/tmN�hr��Gͣ,ν��ff�H�޸�:�#�r���4з�����۹�"�L[���N],�!�I�1VM$|3'�K��~���9�z/b���BP(	��*����_WPth��?�������2V�����D���.� ~��ql �5pZf���9k[��Æ�}��e�8(�(�rעp��?г\u�g�r��'��z���ld��F���Ľ�c�p�p�9>PwH����ޫA�V��u�RS���w]�I�*2�$^f�cqF�P����������K��g��c��{*��v�ik	�g5k*hʳ?�[�Vmr�[���4�6dm� ��G��ݤ�AW�u�.���I,[YY���E�;���P�jЗSK�C�Q(�~�MGba
q�e��Z�j�;*�4�����D����fu�Z�1��N.�2�iy�%s��R���/U��(��kf�����)Sŷ]���k��{Nc蠎!����D�E<5��Lq��ڍ,�#�o ı�F��.>�����`��l5:�MK�Y�}���ҥ������tK����Z�\4���%�����=���~�%M�ιͱ�;�ǅ��lh�=XP�_{����G�W��k����
#�PAq�7B"h�{M<�s�ɳY^�g�����ݙ6eA�H%�c}(D�j��L$�O+�[ĸ#q�Z�F?-�&�`��c瓠"+�_�6e+��%^�q��������wDf��ٯ=wڜg��4��V��%�7�c����53BEط|�t����3���~d�vzݒ1_�h��+�0&����#%��cIz{Z�	/����N�ߊ�QD�<	:�\ �r��k.f���ˡ�n�k��'B��=���[�I�ڳK������iH�h�2r6S5���q��ԐPJY�3�k�?��_�t�y�5��CY�eFZ�`��q39�|��qW���#{2��뭡����M>����P�=bwh����'n5����!�i��Ɣ!O��$y���0����jDJ@{�-CS�Zv�5��,�X��Ia��h?F���f^���6�po��G¹RP}�s,��54-�?㾦%縻�'?���{�cȪA"��^�Z���]>���zh�)m
�\1��!��Qv��hU�W�e������!���p#��{Ѵ�1ah�v��QX�4���V�
��Lǻ;�<ܐD�h9<w�x��ǰA
�i�vor@�����a�J*��A4掌?b��7�����%�>�%������E�u�<����>:0]����=8&@	���'�د�����V�Kפ-����e#^���2
�)���ǝ�RBN������t�J���Yd��N��I7�c_p�h	�
_럵�_!X��"�bԳ��@���	� ��2�T�Nu�Ϳ�j�C�[����]���Y|�3�|��F�#� ���fB*)
s`�Y�IjĭN@_LC�DW�O�նtJ��jo������Ϗz�4زȕc�N�~�b�Ǖ}�u�c��M�A.0=w������L݄@k_��2Mc�-,��@��0!�K�^��Ҙ!�Bk��~�D�u���R�şX���<�U�7�X5�y�j��O�D����O��g�$
��pXk��t�]�g[�ʑ�)������.͐��)З��A�^ʡ�s}�'�-�DN� ��j+.�5��<O�&k��Z���6y3r�L��<���s����x���	��d��{46E��:b��J=ͬ�`%5P`���+`� 7 \�+�n���ki�g��n�´��ʤдV�o�8�l!�s��H�]��z;Av$#q��Џe)�%�;����4����+Q�6]��zH�%���;�m8?˾�j�y)Q��ys��7�1aQ��4W��ӕ��E�R���ŝ� �15ݤ�~�2�