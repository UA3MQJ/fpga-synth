��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+ǚ��.n{Q�̅Z����&�;3j6dED=�Cl���ȸ����8�^+����K�\u��䵌��#���h��f������p�C�R{�`^;:k:	>�@�!y���2D�,���*"Ɯe5���0��ρbL�*�`��V�vX�#
W ��0��o���^J���~#�A��~�.��#������k�h�np�ߗ�"w4�1G8 C�r��gW�e� +�~�nj'%1�f	Fu��#5���4I%�����Foh�s�b�إ�X�Fi���&B%̩�C���8��	�<?��4(V�������ղ���,�dLzeM�T��C�����!�r7�Ж��ڄ{wh3���K�a����X��*��7�8�+�.w|��Mi_�\(��㿖o�E�i�>d� �8��'�x��<�5��Z0�t��f&�/|��{�����TD�0e�8���~�Zf����A�/~���������ٶ���G�� ��d��L����^���骥��v���k�0�vİ�)�X3�̲�f[}�ΧF��?P<č}t绞D�:�����S�K2�?{*�M�}��GV<{d���['4��56xV?�Ћ��+ɥ=��[�
�U�M�uP}��G2Z�M ���C1���Rr�ge4�ח�6M���EJ5���kj�C�i�,�Qq����g��qv{Ǹ?�X����B|��2�l8�zr��c��k;��/���*�N���n��O*f��������}�B�W�g��`H0�eZwn�Z��.)CǓ��_d���_wT'�@8�r\*6����i�
�<D�U�#uW0���m�
`�"��b�@�sII�LS2(���;�և��=g��o�p�\&�
 p�ML���Kk�|wP��Κ����<%�˯�_���t�X����!�BC��-�pL�u*�5٘��O��Gl�p�\Q&O��dE��8s�@�z�n<������g2�H�Sb�$�agm�7J6���W��s��,$R���	!�a���Zp\j�0bZ*���}�7�l�y�
v�g����>U���������wx�or�k� j��S�n�!Rƽ�ډ��1�u�t���x�<��@{�>��ū�sYV��WVⶰ�m>HSړ3Sp�����{rG����|t�R�]_=өrr͗�z�V�*��dF�fX�.B��j2��֊EN�/��uC��܌,�"^�4�3M7.9��>���1�� �z�9�=�$j�{q �I�W�ƾ?��'šoY�1=�o�U$�F����I�c�"��kNki��@���i�C� 9����̍�Rx��\��t��oG���SP�!d`����w����熁W��cd0��阄9q5*��y��7�>���Y� [#��#�@�l�hϼ����JO���Hx�?�a�u����C\>>!`27s��Y_"��\g'MwkL8Øv���{F�Nt!z�����O�Q辫���06���F|BV�D3g� �~#�{�ƴ�D?�j-�"n��[P�$�
�T�В��ٍi�ٝ��_+��f�	J���
�H0i<���E�z��&�k|/�#q��*]5u�Mn��N#O��0-��#n�����vo�!�8�P E]�N������^ʤf�p�?��럢��G�p�Z�b��+6��,�T�_N�Ɠ��A����@h�����DY7�E-���2ѝ�>08td���BU�x���%̔� J��~;w)�+u�&�?<���f�y�G�8 B���}XZy�t�=o9�+[+��������`+�څ7�.X$E�����X��U���i�V�4�;����y��2��"mǋ ?�U@1Zw&H�6!ks�݂c�\)�|��21��g��BU�tZQg)� e!2��/�o۬NA�^� q"/���
������~�q�|�?4*�V�{w������Z�K�j��y_�=����ˌ��o�W.P�G5�M�'rݠ���,��w��<(�|�
xl0u�Q�Ilp�ģ���F&�u�z�"IfO�<iZ6���zZ���o�-��bf@�\�'Ͽ�d��ю�&Y���4w]Հ72�sh��E�,�S[�w���R��I�˒dH��s�x��2i��-��(0obr,��LI�4�(�a]K ��X��C� ƞ����=�&e
����`�ƾiNqؒ�p��̣���
�n�6��M��m��I]r����#/����6]oY�M_-��-?*�r�_p�h�e��z�����K������H���S,
MyA.�.>#�D�=��4h�؟��f��]M��:U��Fw<oh�o#��X�u����s��F�O
�Jc0�L�[�n���v�mI�y>��n���"��)��qB��I �Ҝ�����x
_W� ��ª6���-z�����F��Z�1� p1h�A
�/�}BvKL'ޯ�ޱh�M��ϯ�2G�)U@�PfjQ0(��LB����Y�m���^B��cNd@�i0���b��P����w5ǉ6���&� �U^.����Q�v#1񰼶i������'�)!�O!�3S�����D�|>�곩��O�n7��J��d��!�bK՜H�2��8�ݺ�e�G"Ԑ��*��~�j��]d1���xQ�ǔp�6&�vo�%�'	��&d�./��	����՘�}��=*��l�6N$��o]6A�^��j�ܗ�$hOz~qië-sHvKe7O�E�q���{C��@̼���/)E1���l**���i�G��3S�j��Q/�� �ꟛH�C$���"}��6:x�W��E���8��`�\(s̘
'-sHb�ҷ���5O8�C@�oo���Y�\���.9���)��d}�21e��d���8;*h�űΕ���ΗP�7�������t�FH�����fj\(�a,u-O�8����z�/A�`���1�8�LE��A���{��X�Lꦛ|�8+�mB *Y��C�J�L����+,��8;������z�I2󺂖c%<�0�f�>=�j��I�����lI.=R�
���UС��\����`,o#TS;H=�>����%�WP��2�=����e����ȘE����?b�J�m�
��x��d�[Do�Sy�^`H�*TCkF���ހ���a�Y�&cK� ]s���k�ӰN 9�����~<�1��v�\��C�C&�*l�7�0ӵ���r���|Ǹ\�5�}n���J��k	�d�Gj�ێ�59���\������w�:����Ƌuʏ4H�m�$�ɡ�v���+ay��	� �9��Z��������%��.�͊>jDa�ά��)��k��rH�� sz�����]l�Fq\`SmtNQ�@B�t���b�4�5�>��ӓ����^�f�N�0RK�;�����izF����[5Yͳ�ԐQ|b��'�y;;�9�M��N��j�!P���(i�#���j5�z}IKu�"��{�Ĉ����9Z �M�_C�Ԯ?$�ԕ�k�:���ioI��W�03"�!{c'��#����ڲ�Q	��l��WѩO�B5�W���W��э������Z$Sr�Xu�z����O��5&^�����Sʡ��ȇ,�(�,=����bM+����`�4f�O�/��v��LF�F��w|4(����&]�ǣ�l��1��?u`>m�mK�ȌP��֯2KՔ���Z�T�RJ	p��[�D	{g�u�@�ZO��R5�m�I�8y��4-v��ڄ���p�~H���%���I���W~�솋�\���&Wt�_��߆�i�-΃�^��O�����+�/���A�] ְB���P
=��ؽ�� �WJ·<y��P	�\�_�[!i�� '��ݮ��CV��Vi�<">� ���L��E{�k&���Ӥ�m���ٻ���3ݑ,9�qQ�	�;_AqY�F�1|?9��~�"Ŭ�?G+�e�=@˃>D���'^����_\֌�e�A�qꊸ�'F>;<��+������&�{فy$�M}lAʹQ:3%H�Lp�ޢ?#�el�/���Kk'���$R�9��P^*ZN�-�Ғ	[�ftS>�gtf(CJ�".��ܕ��h�_�k)c�
։~%ם��E̝�T�f;+2�8�O��V^|���ó#04W�����n�L��̍��,�JǏ<sR��.ׯD&"u�A�cJ�=���ºߵJ%�3_�ux;B=o����>+n�t[�aOS'|����I���U��$8y�߭�ܼ�C������Fe\���$��`��-B�P�94>@e�E��hQW*��k��a�в�9S����ɔ��S�.��=#z��,B�Q1`�!Pm#�R	�9�✯�ĘUf+�a8t�DTKk�|q���o��+�M�` �sz�*����Xĉ�]��+��?ږs�\&)]ȶ�SW~Ť�J�D�=�hEG>���ֲƝ+����d�����9SƄF9Ȇo1��p5�+���\Ah�:� ��/�ţ6�1�<<J��&�0�϶�1K��Q������'��=oy�뉶R'X�Ȧ]J?E���OX�"1����H��4�y�g�׈�)2�0Ac��x�i�@N�3��+�j >(�)q���J~B�v+�@v|��Dp���He�>𫃰蹥[P�n��W�-���������S�|��Z�L&�zL�jm��8/���ɷ�)=�`����.p��`fFe�
��aNT2aq'w*�����^�$�^����|��w��0umn�p �\,���nH����[�����I�ҕ�����0*�_���NN��9g�W�-��@�(�3:;�����<StIV�=)��# u'����x��Y�L�*I;���A�	�N���]U�W��Q���pR���!��N�A�M�q�+��iL��$��BP�q�)���Tֱ�s�x%?���>M2J�"k}Zs]��(�[��g$�_:(�$ČɼP��H���oe^���NN��b��g�W,;��z{��4�U�a��U��txK�;i	���O�UҘ�+��%�أ�kPm�4s𣭷kΎ�n>���/�ZO�-�Bx!��ͅ�!!��Pյ�̈́3��3&+^~Ws��O#T��jͧ�P����&��%V[Zo����ͩ[���eѤ�xf����?$�o�P\l���P�O�40q��Ο����G���ne\y�Oυ"���1����J0G�-�3��y����	$�1d���7�I�S�����ѩ�
*tW���zh�3t�T������$�ڙ�Q.��vbr;��zpo��f��J��F%Ȓ�k��w�ٷ��h������آ��h����7I#/�q[ʘX��y#� ��h��I��_�"�|kgo�2S@�EN�]~�d
���v�J���i@��1���k��w�c;���u�d� X��)��w�rao�S�ж7�V�w([�Z�-~]�u1b���$G�s���lf�M7����U��:�/������ҿ[h:�%Ѕ��X	��W�0���(e�U����J�������m ٭�BJ3'��!���1����%�ތk�&���P�À���
Hn�;���?,�\^�pb��:���z+ٽ-��"{�XP �Og.C�{���/�C��CO�Ҳ|�|Ǡ*���e  LE�/�S�gljd�v�͇m@�C�|�ZN������q�M�ɍ��i_��gU�g��
�K��F4������>����KS�WY�\=�9�iHyE�71nbe�Д(�T�e*+K����w<��I7�`0=Du�?Zߒ�<�7�a��'�+��g��V��
:0�r=�O�f=����,+�(O��]���E�qɲ ���6u�����'"ػ�͐��F�i��z���/jZ<V����K�E�����'�E!�ܭ��
�.1�˲O[�K��s_*��p�F6�+�=�EZ6�JYЇJ�?c��#p2˳�K[;���ՄߑD���/P�}e京�[��@?����d��Vw��� ��Td<��_�.KZ����4h��To���F�}����'�����ف�k�;����{0UL.�x��d>kw��5�jB��Mh�r�t^,JI����ۭD] ���ի6H���81��J�b`p�#�U���|�8�W�ݻV�A�D	�1a��)�?S�S�y�~$���G����]=�-����	�-��2��B�!{�v�q�l�(�o����PԲshqY^�ik��<,��X����g�غ����i���;#fn\�{��rh%�)'���T&�D0۶J*�B������W(��-�
��9|��������
v���h������MAlP����z.�3)rv�9|&}�y��|��#d<�L�Z����<!��������.h~]uA�