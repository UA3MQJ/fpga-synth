��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e�=���)C/,��b�IWt�1+����@���d�Mg�d�`�t��_�Ȁ!�0h�JFkJ�S��;�]����w���:��6�����4^�T�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬��\���g�`U<RO�sE�D�6��X,�Z�t�Wdw�%�*��C7l����3.V��|��{�$�H�;�+i����Z�$���p��()g�y]�|�j�4�:�Z"!����X-A�{o��-�Ta����8��I)X�5�:L�\L6�y�]�j�?
������mT�)I��B4V���W޶�[5X"CR^in��)O��/Xew�(g�5l��ϲƥ@Q�h@������4.�u�b8�e�֙�d}�����F��B��^2
����һ�OﶸߑBЮ���q��pه�S�]�;%)Z���97ٮ�6�h�B�5m�* �5^��$ ��Z��\���̴��r�5�W,t]��������>����4`��%Q�����.�r,.d�˛-sbaW�j����/�s>y8���'�Z�`�N��)�I~ɴ�Xi@h��[<�*U߮�lO�Q��ॾ(������,�����Á� ��uJ�O& �re*J��ˈ�O��^Sd}���[8s��/�$2��4S�(\X�2uz�ߧ��5f��V}|W��+s,���t]��(�F����uip������ ��
gR�_X%�5�'T�Ќ��-�Jq�;�s������_&�����r���CY(u�S�,�Y(ٶ�V�<T����O��e+񺌋�YC�7����2��iF���Ct����R�*�z��5�ƨ$��DB��:�~�e!VH&�^�qs�r���"�@��Y}�ӓ��o��s�=.�~J�ׄ����%M���s��a���%����J���qm�Z�������B?:��Y��PDS�	��E@�g]S�/?
�"��H��t��K���x�S�h����gceP�cy�j!��PP��"*�B-^���n�nR�����b��
=%��\�s�V?ñ���֭�
a��L*7�Հ��Cҁ�5�4&��ZGV"=v�j말ЬT	���1+�x��׈ߗ��+����ڴ.~iA����`#��e/�ī�z�d��r��B� ���3�
p��2+?Y_��rg�P�p�9�A��x�ʫx�2��9�����K��K8�
a�K���h�#!�����\F'��:uҘ��/�г�/���{��%�P��q>�w��r�[q&r�FA�ga�Z�CҰu�֝�k'w�2s,���Ҳh7�KP��1{P��3�-8�GG A�om��!o�ζ�e>��߫��}61<,������`��쪬}z����!�ߡ�8�(���*�m��D��h��%�]�w�`��2�m�Q� e�oD4c�FZ$�$�}u.(��?s�B"�*=*����$U���Q�m�6��'��8�d�p�̼���7�'d.��@�N�WJ~a�PO��^t�XG �b�Ke!��gL뭐�Q�'YYXCb�H�}rJrm��-�/b�Y�� ���Ȝa*,�oS����f�p�hH��*���=��ۮ�$�̮W>ζʁ�\2gZ����[���r鉡�����tO�Ǒz  ԄB����Da.Y�ٖFk��{�Z>�x���h{GbI)��Er���[J��QGW^!4���B��NN��i{������7{&M�2O�Xq.� ��|� )����

I�J�'q&�+�#�r�p�gM�hܼ��KU ����d}jXx�C�o���!���1;:l�]{LC_V�lc(�����Z���1u��)�&!�A�6(�B�a��æ��������a�Ə@"Gto�2�A�m�p���I)_g1In�*�l�ԞOwpiƉ�b�������I'B[rP�ң�D�-k6gL�Vc�����d���ĚO?��*G�f�{�d�U��n,
B�1�b�Ja�}� �	��Pꅔ;^\��w���]$�]3�}����P-	.���ݥ�%�n�����,�j
F,�qjvN�[+$��X� &����)ip����+�.��>�	�iˁ��[�d���1��d�D� fq8�Ϙh��<��In�&}��.x��EX�x����ժ|~��U*�T�;�3���<�N{�]��e5�w��������4ۿ��|$/(�H�$��G^�y�Ʉaq������q(Z�C���0�L
+:���K�^^���$���oEK4K�y�m��l�O��{`����~�'p?tx�}`�/{�JK.7��F��]���2а��An�-)R6[�\C��L4K�;ga4�[�f�P����`&#����h��wI��x�
��<���� X�0b��Lq��7n?�=�/Z�l����gm�iJ�Qz��3��з�Z[ȡ,'��y�(��QnL	����]���w޽QX�ֲ��dpu���9���\��φ��2�j��(��9�r����� f��5�B/�����{�����9�Lf4\���#��kś�x�"�s�vџa�|�K�g���`����X��?%r�*� ��[��fVC��ů_�B�D�;�.���̋'޲qђiy��D��U1��L�3�Ҟk�]��s�`��ه��`B\@i����]/�'�Ņ�7�e�ђ�%��n|Z=av�PL��"i�Ⱦ�V��d"T�b@^hZEd�\��e�������~z�&;�U��0.��9m[�k���`�&�(i��3bif��tP����^~+�iYe���X��
U���Ġdz�t�9ʬb�_*���'�	.�q�)A� ��Ɨ'�:�Xʴ�����D	�3�G�o�=c.��j�&	W'�L!�a	d>�͞�:j�&�QX]������:Z�oK;ܕ��u�	���<��,��r8$�n�����T��*���WҊN�)!n�`5���n[���ߎs���L(��.Oۀ{X4�D�2Kd��ŏ�Sd.�f�����^>�"���J��mt��
�����cV457�=HA�z(��o=ty¬��7�����V��CtF���t��T.߷��c�\&��W��m��p��(,���р�+��2=�Er5I�l%~W~&섣�� �Ts����^�0��ͧ���ډ'L]8%N	��N$�_Ue��5��w`���&�T��G���_���`��vM>ƝH[�$ѓe�o�OT�y�d��>�5�i*g"���l���� �iin��q���~
���~S�'<�Ӝ�`M![CIA������|l����V�T�ftY�w4�iܖwiܵ���-�	�J# YyKV���Q���f��l� z�Z�5�]o9��޵�V�{���Jƒ-K.	��������<���	��ϕ�,4}���H� �M�)�[|1�J
z*�it5��o�_�h��d����"ǧ�Xc�Q�h��v��9�����B268��+a���FU��۳��ѿ���U��SM��3�g<��1����ܮ6gj��yf�`�r=	4+@�>{�Bcb:�I�vob��Gp7��pX!����jaZAe,�u����2f�6�M(
Q�Z�ϕ�޾��t<�e��Z���С��v�SPD��B�w�O�|tx�cP'ލm�#��~�)�Lm�V�V3L�;�q�hڥ�~~դ-Jx�omgH�x/n���>�<��Nds�"����yf��DH��ƨ�!�����~�M�.�`������2����~*�GB��������jrm􍮀l�
�Ã����p�<U���)� H�j0�Oj����rM����Ec#�U%���B��w�����QM��
� M&�A�	�� 7���5��YRnF��B�������~�-���C�/|�� 
u��k7&bkK�+��%f_{�[<=P�2d}�C�p'(ߋ�(��)�M��B�n,X�=쳕��5}�����}*h�<���ll�e}ظK��Ie]�o㰌&w�ھ�Ģk�S�3���7���nHr��ɛ��^P�ъ�v������z�M��� �L>dܯ�/8�B�Q�}�G%0l��i�_웻쳏�l��l�{Hi��]݅�nXi�M��w�S&�-�_�iHd�y�ڲ~5m�����9�4&����ܳջ]�E�/�	�M�8��Hp4(�Yk��?y��ʣ!CBM��'�=�8��V)�ǌ��m�斮̍~�+*�hf_�
�/��p�yyӝ��ib��&��nw"���t����/Ͼ'���x�J��^��AI�VU�5_�H��n����r�I���>\�E ��q�o��p�K�(C�y%�W����Ғu��JQ�D ~�$�z�۱>9��(�C_�0Ca�L!ʐ��GZA�~���=�����\��n��d�@�#�+�C 2"�@$�\�?3���!�w��1�>ԑ����Enc��OT�e���Z��FU+����y#�/|=�W�
,��'Wa^Ѷ�4w��Q��l�Q����R]��.)�d��rL��#�Ym��@WW[!]��Zi2��Ȧ�,>J�蜒��1'�~X�,ʷr�s�0��_O P���t��2o���a�a��'�( RP�E�\\Ži�_�[h��H6|/s�*����3i�	ᨨ�p6��PUIo&�i�َ���w 5�k£��{=��߳�&���n\�C8K�"��|�@:X%$#lD�c*�ou�w9���_H+�Hڙ?u%�4*)��·P��xXp��h�=�E6�s����Ի�X�MKэ����x쬜P)��ļ��Q�2���a;�U%��c"	Ԍ̶
�^�꫶�����NjG�F¡���Z=�
�� ��G�r��X�^LT��o�h����~KW�l\���o�)P+>�K#�l�L�M}�ֻ�[� �y�2-��ɪ�mX/[��i�
��/�y:M�iiO��_�Ӯ�/�8'%V���C�%����b@wҴ~�l��d+m9��	�v9���H���T].�bow�����O�g�#{�+r�H��$X4NR��w�!�YmP��u�� �w	,���.�a	tf;T��-�̶�͋c�[�b8��ѻ[e�ȿO�O	.�>;�-�1��b�~�I8&2�7��	�H�Wu��}E��>�� "@SUiS�5c<u�<[A����L9j�|9[�mGZ������S�3���CE3��@�,*`�c9l].T�jnHWeA@d�H@� �ecG3v���rk��n�JY��UP���r��S����-�^���������!��ʯ%<���=�S�ё鏭���oK5�����ʼ��(�F�J�����V�����D�S�ndsp�h� +K7��,�)+��n*{1�E���/�}^(YL��ݘYb#[�z|<��	W�8~���N�_ƏZ����I�	���0v��}�%���/b��0Q�I�gjMI���>F�D�im�����f�� ����+��/w$F"���7z$@�SJ��;��� �Y8�RU����R�T����K(�4\*����W��坱-�o��	����1,+\]RP�i%˿�v@^�� �csB�vNn���#��
�V�����f��>��n�N�ҋn��r���G�\10;�r�R�a�s]`M��K����$q����o�'4YOː|v,ҁz�Ҷ�Z�Q"��<D�0�F����Ʈ�25�ȇ����Y炳��UMG8X+�y4���#@F���/�B��$} �T�3�F�j
b�<����;}���j]�ESP���L��O��B��vc��:��&�M���E�K6�u9��~<�u���F忘@5%�#MT�	�3�TA8|,�'z���oLG���ϭ� DM�4����~T�Ѣ�6����ک\��V�@iV�؂�M�����M���0W1�(M��匤:�;�`U	+ː�Tl�ancX�E�/ C'��PX��oqoxT�U���;h���M�k�Ӑ�U!�
*f�8�+26�Cbl'��U�e��9�TN���ٹ�ڛm�з��PBZJ(Vj<�����/\�_��]8a�8ɒ���U�f}L�9﹵aX�S)j�w�b��o���Ǒ:h#Ͷ���h���w�$��+6����g���� ���ʹ��qzS40wg�>�{S\`6\���p\��:ޕ<np]����C��M%��od��6&��jF��5���%�w�;��_��e}��̄�����g����kM�� �u��o7Z�8�̣c�:�o�0�kV�1���l֪K�:YL�Z��	��]��Lj��2+m��n�q�)U���c��4�[ٹ��s{�|��PdМ�z7�D/7�(ly˺���uq�h���7�`��J �8�<��C��s��N��L�ԅ���E�Q|��D�����-_�=Êy��m˿C����n�p	�;��+�|����Om��� ���J\�L�͇��6`"��f��H)��e������L<�Y�X���҅�I`��c�A��H�.4
��$]U�p��;���Eԥg��$Z��o�gv��������i��-�:�R�EbF{>Q+Y��*"���vf(ה�$%Z���g8��J����O�� �GRvⷯ��M��v߶�V)�Ƣ�)���A+�9CF����(��6)����n'��F�	H�������x@�@v]�m��^�_�e>X�m��oS[�"�a�������C�e�Y?>Z�<wq���e����F<g^��<�p�a�dR�az�����Qϖ�D�)��p�zw�Z47[̳�]`΃���w"I�4، �tH�C *Ê͑=~��b�6w��7H�,�K%ް�]!�y_S��?��crmcF���f� �v�͍br����X�8��I�Ig6��j�ޟwx�4KvI�!~U�R(ϗ�H����lu5p9����u�T�b>�X�����3�~V�G��;�Q��~>H>(�n0ƅ�&\���6�q
먥_ȿ�b��`҄��=nG0���%��z��'PXF��5MXqJ��k 1Ŭj�����L�b�*�mOرꚴrP�T`溺n�s�1�-��[����K7Mvh
V�Z!>�*S)5���<?mivLA�s���gj>�j.�6{Q�G%.'�T,#�@@Ǝ;Lh�항M0e�������ћ��?�n��c&�%|yJ�-�(����Tl;78�%b��m�aY��K߶k�ζ�0/ݿmo��������������1��Y��K�q����u�}��a��';:����W(����)�a�������M㈌ʻ�y/�45��)�s1�SyZ�W�LQL[�+;�"7�V�H�ۖ;��_��lP����N���
,�w�N�?'��z�	�������~Ǳ�}��1����/w�)�7R��j��ʺ]C�v?�B�A�з�I"��A?��c6:�{�u�H�_�ؚ2e�I̚�摘��{�m�!�� �����Q�&�K)f8�����0���,EЧ������׮<��IӃ��Ζ6(�kI9�DoڲI�xP/�g|�x!���*_mC=�c��s��ĵps9��X�o��*��j����]� ��/�����XH+&)�F�����4�x�F��x3.GLL�V�S���la[)���N�y#�m�RFv��*�(����uv�������F?.,���#},��d��E�'#�������R��tk����x-���Ծ&gR#	 gA��t4��P®�ܢbZ�B�N�ٗ��R��f6g�)q�&�қ��Ĳ�����vLw��X洓�?�,X�d��u�ݛɔ~���l�h�=�h�����MN0�ZY�fa�q
�؋ɵ�v�;�B��C��9�~�"a�-�Ww&^���_$y�˦��)O��M�FX�ܑo,y�ڽJ5_yI�iq�*_j�@����$�J�ہ���@7���ߙe�av�*eE-W"�e0��'�R!�_��HEr{&J����j>2N��B�	,Y~0�����ϊ�ur�k�Q�c�/��B��y� �_�꧎�}��Z}��dǽ�<�3bBZh"l��ƕ���R_��`����=οHL�⁒&(/���C%c��
�Dg�7\8S��y�#3�G�]�tE�,!p��jʡ��44m'zք
�囡��ص|o�0��,���y�!�C���1�Jn�By������01uGP����}ח��Vv>^�1�wL��b��� �,�x
��j��y�7�z:�����H����y�u1�	ɼu"k�+j!���g�ؠZ��O���:ы���>Uy��ߝ���?��G̑�
,�!����iMk�ِ ��srD���+F���I̮I�!g���������j��5��0Ad~U;Tj�������mq<�r�/,��7�B+ kW�Z
Ώ��h�����׉XL@������Ή���\eK⭋#���'wJ��IE�q�@��9Ŷ�X��J,V�U[�!����j��L
M/����*D.���nH5CwP�4$y#͋$���d�T���T=�낮����+�U	�t,��,���zT^�$�%���7�Y�!u�%�UNh�K�ND=�%D� �r�xCj�k_DT��Yu�5�t�Uˊ�9�M|��|���� �Q�NC�pq��:� 4�$�ۂ��\�:��0̡jC��ڋm�Ơ�+�])+��%�b��?m�\A�f��%ۗ���,G���2dԂȥ�9�����}�VU�����a,�`��H��W��n���y �:S��=acH���뗢�	V w0�˂�\�5��f�E����$��Nl�ڸ1X/��fz��4Mdtn3�����V���� 
�ϕV��z&�ŉ��3%�\?ڏ6�^9ؤ2�_���r�|px�$*s9u�w<$�=h�H�~PRi���� l��4����fn��0�d������TI3��z�N$����m��,��#�Uw��Ƭ۩���(��~�YLq��⦋�'�Uj��?���;_o��6,瞦�g2-�(�u������
�Q2�[�2wn���Qw�v0KiPF1�GZwӡ�12�ݓ��k+���V���R���T dT�W�N����>l,�Uw~�H�in�z���'�*ǘ��F@���1�)O���8����G2v�;�uO��;޺��1A��0�/�qU���=d���J��*�G��K<f�_�·RsF�����|�b�-��_�B������ ��[ۮ�H��=�wL6F�=KՔ�?I����������)n�r�^k�R�7�QB����~:�#��=I�a����і�m�8
���6�tO*(����h�g)74f9�a�+��+R����l��F�:W�rI��64�-%Hdn.�:v�s%�X�a���<E����t�D5f�4��v�OƨFB�pg�0����a
&�J�xZm���L�b
�1^q7LI%!�f��HL/^^�tIh}!��C���1�ȩ�|�c�zG�`�\��:����ʵB��0��1G�f�%�����/z�����d���IVK�!be�0��'���~�z�P�s	c�X����;�W榉�^;�!�X�����/ݽ+̆}p�r���]�-ڷ��=`t1��Z��h'П����'�;�8����Z^�OO��v��"��J�+v�V�����]��M�����̸�T��dӋ*��i֭]���U�Ž`R3X!�
���Q�ܨ��|�@3�f���}ܰ�.��QvLm2
�ݾ����i���̉��<\�[�Pr�PYx�Aү�o{`H�~���8k����!�h���wGD��5�@z�H�3��=ukc����0Q��,�vI���D�Ԋ���MG�k�4�tEPb	��B�b;3�ԡL �޿���"��vat滥��A��><����\8G|S"ܬ<�UH���犀^XI���hIڸ�i�9���U�7��"�8���1�a���w��j��%��4��u���D�4��'#��R�A�����9|�� ��"F��Ш�8oh�.��!
�LDaِ@8P&8���萉9���%~
 /�3�r�A���3v\1ƌb�f!V&�!P�����^W��@���Q��|��k�WK)�#�1��s�xQ���l�)k�ʰ�wRv�o�����]��2Re��r*���ث8�U�� t?LX���4�/@�
��U5���>�z{�p�]�'P߾�o7d�u���t�+
k����w����6���B��������}��U��|�@�&�Б�e�oȬ���(X��1Ix��#��Q�J-��SK.�v�07|�C��v�.�f���4��}/�0Yڐ��SW|�b0����5���*<9�gu^�x�|��zO���Y-�3,R�]��<�-2������g���(�9eb�/2K�Bfa�Aw�}�z�����΂���m�˭#�e�a��@u��"!���ݥ��ekmu�F�n�Rh�oЍ�P���:���bo)�
,���}��������s�� s
�DC[��7]�hM������EJ��@���D��/��v��Lß�ˏ�����f_1׉}�>o���j�((�j�cn���0�W�8�.����2�3͗=���V?�Q�����s�-������7㭭+�kT��W�E��YO'�_��
z~`�������3)��t{�ue�,��_d�x+���*-Ёq�|�S�
 �_Q�},�*�䁐h�k�gZ%`���D��w���Cx�y��N��z�d�1Mb���S�g�� ���Ҹa8������dMz�4ƫ��ޮR>L���0��Ԡ��3 �\�@��$d��9�ۛ%\oߎjζ"��Ǫ������51RboK���^b�����#���X��Q/�걁m�����˿�z����p!P��(�!_"z����5k�=9i|�޼&7�D��<�'�
����lm"Tk������|!���eZFO.�mgq[	��H�EZ,p/����swϋ�㬓���3��V1��4�9���e�-��Б\͵��4c����lh����0�ƗZ�� �/�ڹs��$x�Pm���W��f��gܭ��;
T"��J��[Mz�e~Cd����^ط���r�܈Ϙ�'-¨-53y x�<x�*g��ɶ�p�}�����L�M\�K�@�\mb�k��Rc�(�ѶNڪş�u��kI����\��.��;���n�k�{�b��i�UK�D�u��F�0�3�R��"�M%_�i�T��_��Sӯ��p����M8b���t���io��Z;�Ы �f��˧��$�� ������[� +�b�Bn���\����)��g�;�U���J�{�qW;��B��������4���J���v�B���F�������HM��ҙ��g�V�0��)�Q���h�bf�A����PA=ȭ~��~�6�=Ǚ�����
���c�a*�<�2�/�JyJt8L��M�0�ԋ�TL'�>���W~�掫@�h$V��hF����4(��6�W� ��gJ+ �y��$
�a��`�B�..n�� 𯪌� �?�Oظ�G�Ϛ�U,W�3������ p�3Vo�!�l�9c�����m	����I�"���M�o�0����!"���%�H�[�]�Ӏ!�,�4�S�家��*�-���k�Nt�.�$R�n��ݻ�@�q��R��o��p��]��}H�	��������� _����9�X�Pv]��c^�Ϻ�"܏��l�VT8q��}��	�\a��$ʻq ϕ]���T�^�C��wT�>ʏ{K��v��0D��5}���\g~:���P�O�%��H����b�l;���D��w+��{��.@� �Q	sQM�'`#������R���괲נS���Hp�P�P��] Yyl��w��Ǭ�n69�L4>�ժ�9B�ݗ�3�!�ڲ���'��S����AU� ���t���L/�!�����ԛ�p��Hg��lT�K����X<����I��Y�c�>��.�d)U���2�q*Ӱ��,@L�`2�h�RϠ�9��h�ka�0��I_և@���. ����+"��G�fJ���jWL,@�*$�7R:���8p�^ܴEU�+�����D�ї�W�����Vh��[�T Y(��a�;��b�ĵ7�9v���!�����9]���1|R��!/�s���}6����70?�@�z����0 !�ƴy��C����h���I͢6��k��}�T;�(���X�N�TM���+؄���_D���f=���
���2��: �} k?6T�veI�ŏo��#Ƶt<�Ǩ?�A5����j�B����A!���滶D����7�s��&��b#�z;��ʅ�;����Z㆚��=��@4:;
'�)�+�,�����bB��b��6��[1���VV	j��=�#E6�$��� [�3��]�C-F�|��փ"/A�tCV�6�S�a���y2���]���#}��u<]c���,L�A�3�5A��S�]�U^KMp�B���P,�/?�X/��/�Z�L�%�I�!B���P
�rn�3�>[;S,����l�QO���@~�|0j�nf��m_���|����w&ؤ���G@�R�%�e��b�;ع�y,�d܍�BD�0Y����u������e9