module lin2exp_t(data_in, data_out);

input wire [6:0] data_in;
output wire [31:0] data_out;

assign data_out = 
				(data_in == 7'd00) ?  14'd07540 : 
				(data_in == 7'd01) ?  14'd07110 : 
				(data_in == 7'd02) ?  14'd06704 : 
				(data_in == 7'd03) ?  14'd06321 : 
				(data_in == 7'd04) ?  14'd05959 : 
				(data_in == 7'd05) ?  14'd05619 : 
				(data_in == 7'd06) ?  14'd05298 : 
				(data_in == 7'd07) ?  14'd04995 : 
				(data_in == 7'd08) ?  14'd04710 : 
				(data_in == 7'd09) ?  14'd04441 : 
				(data_in == 7'd010) ?  14'd04187 : 
				(data_in == 7'd011) ?  14'd03948 : 
				(data_in == 7'd012) ?  14'd03722 : 
				(data_in == 7'd013) ?  14'd03510 : 
				(data_in == 7'd014) ?  14'd03309 : 
				(data_in == 7'd015) ?  14'd03120 : 
				(data_in == 7'd016) ?  14'd02942 : 
				(data_in == 7'd017) ?  14'd02774 : 
				(data_in == 7'd018) ?  14'd02615 : 
				(data_in == 7'd019) ?  14'd02466 : 
				(data_in == 7'd020) ?  14'd02325 : 
				(data_in == 7'd021) ?  14'd02192 : 
				(data_in == 7'd022) ?  14'd02067 : 
				(data_in == 7'd023) ?  14'd01949 : 
				(data_in == 7'd024) ?  14'd01838 : 
				(data_in == 7'd025) ?  14'd01733 : 
				(data_in == 7'd026) ?  14'd01634 : 
				(data_in == 7'd027) ?  14'd01540 : 
				(data_in == 7'd028) ?  14'd01452 : 
				(data_in == 7'd029) ?  14'd01369 : 
				(data_in == 7'd030) ?  14'd01291 : 
				(data_in == 7'd031) ?  14'd01217 : 
				(data_in == 7'd032) ?  14'd01148 : 
				(data_in == 7'd033) ?  14'd01082 : 
				(data_in == 7'd034) ?  14'd01020 : 
				(data_in == 7'd035) ?  14'd0962 : 
				(data_in == 7'd036) ?  14'd0907 : 
				(data_in == 7'd037) ?  14'd0855 : 
				(data_in == 7'd038) ?  14'd0807 : 
				(data_in == 7'd039) ?  14'd0760 : 
				(data_in == 7'd040) ?  14'd0717 : 
				(data_in == 7'd041) ?  14'd0676 : 
				(data_in == 7'd042) ?  14'd0637 : 
				(data_in == 7'd043) ?  14'd0601 : 
				(data_in == 7'd044) ?  14'd0567 : 
				(data_in == 7'd045) ?  14'd0534 : 
				(data_in == 7'd046) ?  14'd0504 : 
				(data_in == 7'd047) ?  14'd0475 : 
				(data_in == 7'd048) ?  14'd0448 : 
				(data_in == 7'd049) ?  14'd0422 : 
				(data_in == 7'd050) ?  14'd0398 : 
				(data_in == 7'd051) ?  14'd0375 : 
				(data_in == 7'd052) ?  14'd0354 : 
				(data_in == 7'd053) ?  14'd0334 : 
				(data_in == 7'd054) ?  14'd0315 : 
				(data_in == 7'd055) ?  14'd0297 : 
				(data_in == 7'd056) ?  14'd0280 : 
				(data_in == 7'd057) ?  14'd0264 : 
				(data_in == 7'd058) ?  14'd0249 : 
				(data_in == 7'd059) ?  14'd0234 : 
				(data_in == 7'd060) ?  14'd0221 : 
				(data_in == 7'd061) ?  14'd0208 : 
				(data_in == 7'd062) ?  14'd0197 : 
				(data_in == 7'd063) ?  14'd0185 : 
				(data_in == 7'd064) ?  14'd0175 : 
				(data_in == 7'd065) ?  14'd0165 : 
				(data_in == 7'd066) ?  14'd0155 : 
				(data_in == 7'd067) ?  14'd0146 : 
				(data_in == 7'd068) ?  14'd0138 : 
				(data_in == 7'd069) ?  14'd0130 : 
				(data_in == 7'd070) ?  14'd0123 : 
				(data_in == 7'd071) ?  14'd0116 : 
				(data_in == 7'd072) ?  14'd0109 : 
				(data_in == 7'd073) ?  14'd0103 : 
				(data_in == 7'd074) ?  14'd097 : 
				(data_in == 7'd075) ?  14'd091 : 
				(data_in == 7'd076) ?  14'd086 : 
				(data_in == 7'd077) ?  14'd081 : 
				(data_in == 7'd078) ?  14'd077 : 
				(data_in == 7'd079) ?  14'd072 : 
				(data_in == 7'd080) ?  14'd068 : 
				(data_in == 7'd081) ?  14'd064 : 
				(data_in == 7'd082) ?  14'd061 : 
				(data_in == 7'd083) ?  14'd057 : 
				(data_in == 7'd084) ?  14'd054 : 
				(data_in == 7'd085) ?  14'd051 : 
				(data_in == 7'd086) ?  14'd048 : 
				(data_in == 7'd087) ?  14'd045 : 
				(data_in == 7'd088) ?  14'd043 : 
				(data_in == 7'd089) ?  14'd040 : 
				(data_in == 7'd090) ?  14'd038 : 
				(data_in == 7'd091) ?  14'd036 : 
				(data_in == 7'd092) ?  14'd034 : 
				(data_in == 7'd093) ?  14'd032 : 
				(data_in == 7'd094) ?  14'd030 : 
				(data_in == 7'd095) ?  14'd028 : 
				(data_in == 7'd096) ?  14'd027 : 
				(data_in == 7'd097) ?  14'd025 : 
				(data_in == 7'd098) ?  14'd024 : 
				(data_in == 7'd099) ?  14'd022 : 
				(data_in == 7'd0100) ?  14'd021 : 
				(data_in == 7'd0101) ?  14'd020 : 
				(data_in == 7'd0102) ?  14'd019 : 
				(data_in == 7'd0103) ?  14'd018 : 
				(data_in == 7'd0104) ?  14'd017 : 
				(data_in == 7'd0105) ?  14'd016 : 
				(data_in == 7'd0106) ?  14'd015 : 
				(data_in == 7'd0107) ?  14'd014 : 
				(data_in == 7'd0108) ?  14'd013 : 
				(data_in == 7'd0109) ?  14'd012 : 
				(data_in == 7'd0110) ?  14'd012 : 
				(data_in == 7'd0111) ?  14'd011 : 
				(data_in == 7'd0112) ?  14'd010 : 
				(data_in == 7'd0113) ?  14'd010 : 
				(data_in == 7'd0114) ?  14'd09 : 
				(data_in == 7'd0115) ?  14'd09 : 
				(data_in == 7'd0116) ?  14'd08 : 
				(data_in == 7'd0117) ?  14'd08 : 
				(data_in == 7'd0118) ?  14'd07 : 
				(data_in == 7'd0119) ?  14'd07 : 
				(data_in == 7'd0120) ?  14'd06 : 
				(data_in == 7'd0121) ?  14'd06 : 
				(data_in == 7'd0122) ?  14'd06 : 
				(data_in == 7'd0123) ?  14'd05 : 
				(data_in == 7'd0124) ?  14'd05 : 
				(data_in == 7'd0125) ?  14'd05 : 
				(data_in == 7'd0126) ?  14'd05 : 
				(data_in == 7'd0127) ?  14'd04 : 15'd0 ;
									 
endmodule
