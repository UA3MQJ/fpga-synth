��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�l�U0>�����զ�@��������L�3X��ɸn���'A��U0��f��݄ �.M������ZI�>Hz�����Q�C��ׂ����!l
��W6*��۶��r��6�3�\�^ף/z�س�����鵉�˞CV�MC��	��FKX()��fb��m�cVF7��=�#T�'�[QwB�/A죢,�D1�I�f�;a��H:W?FCP�C˫�@��"��o�t��8���,��4�`���c��1S�р���n�*T}�ΛnY�ptX�ͮ�� ��r���(��|W�=��H|��ǐ�=��Ƙ%�|�&��&
�$+��~7�1 >'F2��`+P F��o���`x	H���s��@�=븈L����٭J!�+F�0��Lko�<�ѯ_������-7���蕹/�sD�,$��s3�q\ဩ��*�6��ۄ�벱�m~}u>�U"�%,��l�)_G(/vZ�E݃�J,i)�k����>E _�o�+M�(�{���K��������_ĥ�Q�nYk�N�un4/W�G��$�s���5�s;�s��<�VL> $�9^Qw����Wh����}R}7A�����^D���9$g�ONoY��0��ۯ��64L���LҔ\92"����|�6~:e�/=ȇ��E)�u8�!�\�?��@�OYL�;r��=�͸�E��N�C^�H��d�MiY��q�#�2S�{5@m �&,����N�0����*�Z���̙�FC8]��2ƭ���o�*���5a���_`�8��̣%g;��mre��0��H�<��w�Hl�D+�*ku �C�F�%C+��ewD�ӫ�b��z�a���28�b1
F�z��f�T3�%�uP�(��_�C
�O�p�XWoΨ�4���^���v�L�@(��H ��$n��:*���wGe4f{���f� ����XT��'G���DU}�<�.�Ap��/sҎ��7��������הb֜i�S��u��Z����!��u�w���2Ae�e���8k��_U���yf���6i��U�����xd�Od-�/��<�K�(�(�������Ew0���o�v�e\���ڑ�5���(���zywE�&^%�Hb��T��2�;� ��w�.A�Sy@g����>��'U�y�$�+3�bv�˘��$�Ry�g���j���!^����#63���`2�n�����*���k߼��{r?3J���.1�6�a�8���򋻻�&��#qv�A�Ǉ�05�Il���ڕ�e�-W�=����l���r�����YӰ��MEڃ�8����v��ȵV��Q�u�W�;#k������
aL��r���C�#���(�[�l�F`�F��csd� +ȵ6�)����N�=�f�W�Eщ޾��[ޟ�	���	eN�{_'vse�W���%(��A�4{�a�
n����P�uEp��M��'��H�s_����4->�;��Uү�@^TVk�f��������	�)��jeC�Ȓ�w���X_�����Õ5v|Y�z�U}*x�@_�ޡ�@Zl�q����6�(`���䙰���_3�`��A94�pTfa�Jfi����V
q"k��hI��u��2Ls��;jD���&���43.����d:�ɫ�l����p&$9H-1�8�9�=�$,�~��zL�d9�P�V�'�'Ʃ��B#՝�)a���i�pK8螦��h�3��Q�T�rf�l}�%C�ȩ�*�謋G���RK�6�w���-�8�E'�q��v@�=|q��dM�ZZ0�|k��s�HP���mjZP�g��ڦ�=�7����W�rv�N��Эp�	��C�ry^�<��H�;�bI�4�#����\Y��v�Vqǵ7����?����A�W�ރ0��M��� �_nr�����~�X�2x-�H��E)C���i���� �����*��h;����_R�&= �ʫ4�n����Q�x$$�5>��K� 﨤r�E�g/%��5�J�j��U��^4ݼ}obz!�����UeY_M���SM)UZg���"��M�l�i3���옊F֡�u;��ћ"��1o�����л�=�B���}�R�UI�D�]LE/F��_	��~7��΋�ȉ�8�����i��W6���7��s|AŤ+�G�|�� �Z���n�dj{�w�!����8c㖾� ���[�hy4�X¯�ry2�|$�r/��i̋��ò�o���&�Ťh	����Z���{ڔ��
�J�˔I^<�u�i���^���n�T�FJl[��#f�3L$�#��C��|�RZ�͓�Yz|Wm�y�bM; ��E�"��{��K��N�L�YX�>�$O-�y^�|�� ,���Zv1�[��,foX$���B��k|l�m�#�"{��r�V�{HJ��+�*om��׿bI��|O�)!���ԋ��S<�A<�� ��ףA%�~L���G�����ãJ�]qͿԫhL̱Ǩ�Mÿ�>3_5&�ػ��?3e�5>xF�qnf�ix�ξ���b�zxs�t���eE�@�-��1Z��=ۓ��i�K��{���>�HDnV=���H��sg��SD��Z�K�#�"H��;��< �t�	���/'��Ra=.�y��Ĭ�� �3JaR��J�Ѱ�l�i��n-�U"��\�*��Pb��S�
ю���� N�Y��J��RV,Bd^�c3��	�$�1�A&�p�^}r�m(��#z�i��>lKjn!���+�[1�ٛ�8�u��QL�nq����A���U�~L�,0�Ȝg�]��w0Ƃ+�Чy8N���w�M���	,k�wUՆ����/
M ��ڰFv�J��ǫä�m�X'�n�vD���f��$�1�'�ǈ�����|ܪ&6����h#���2�3���;����D(��x����_Q�>,e6���L��`���q�(���J�j�͑1~�	�l-���\�TZW��k�Z��L
 ����;Ff)x-?I�� C�z�1fI!����ni��H���+�
�4�p�9;��&�1����M>|U���kC�z����N�D�4k�?�ĬS����Z����K�a��vq*����e��eʹ��2ܪ�f�$�A4���D���D�D�,�p�s@�e���Y%c��@�Z`�?�\�¿����M�/�i)և�=hΟ����$ӑ�;��F&Ǆ+^#r���I�׺]}�Gv'���MmȮ5��i���,Ѷ�y�J�R��k���s���w����I�#]?��N�����~$k}�@������=`��������<�@9�cf��L��1Pu`i�x���N �+�F��x#$9Lւ��L�ģf6��N�=/;0e�ˤ�_3��^���	'�y�V4���s��f�egP�*� �n�l����W�[���N;=�!$��� vp��Y�k��!X����������m��D��`���"�s�2��:FwCs���ㅎߥ��u[���y&dݽ�Y6e�%��5� ��t�kt�(F;��g�1�J���ǽ����m���$����f��n
51#��f�}Ơs!���C �f���t#K�T܍����Β���?J�P��Ɓ�l0�^?�� �i�?���+y�?��ߠD8YþÇ�JV�^H�s��4�g������8(��m�
�'h�퇿�ɀ>2��8�`�>!���޲3@��.Zx�z�ȋط���E�+�XA��2r��f�¹�rΞL��yuL���9�e\��8��Ͽ��W�a���}0�3F!�GP�[#�1=���k�]Ҋx��ݑ��W��,�ۘ��"��t֐�ye�C������&4���¿����63|����4�ˍI�[�H떺�[2�Q�F�<�x[�A�8A{�����-�>��E�ʗژF�k^y�׻�m[ў��M��J惷qO��.Qub���Iu�%��]i7ᒗ��lj�H�as��6��o0/��\�8[|8m�U/�tg+�f��b�╾|��DH�b�$�AM����]v��k�P�	|'�P�$���+9,��� �ݑ��v���o�����͋`XWhu���X
f��'T���N^�g$
)�l�>�����w�+M�0ݪ<���z���-D?8��u�\�ͪ��į�
��"&ɴO�ׁ)@��?�HM�/MZ�X�T�>�($��.�´&}[���v�x����&l�I��4�AZ����/����(2i��P��`UX�M#v��[I3���	P�dX�p�eP�&ښ��E(��h���1�C<,�X��o����pǙ9�uXD�`��w�2��ԓ� =�?ĭ��4��������W2��:Y��x�1�D�Q֚Jf��@������?�&��N�Z���#��PH$<�6�_��[��fG�< K�ď�� B�e���gA'���PEH�]j���yv�������`��A������"	 ^���70%X���y����܅R�5K��RV	�Yx���'빧��px��HT#�]ձ�9^��+o;���_�&���=�p�,0���뻞c��%���\"�*��!��_�O���#K��0i��rg���.E5nH")�Fp�myH�HO|2��C�D�spU7��W��#zB����WG<�<0�&��SCpat:x��Ԕ���ۂ��@�������m$�XRZ���e,Ԉ&W��?��@�嚮F�܁"(��H���F��<�/N�Q<^h3�0��Rwyg�p0q7�1r,�_Q�Heݦ;zS��G �5a��lF\�d�aI?���ҁ�:�y �";)4``���y0�^��Q>��.�}N(M��v>�Fױ���T�$"�v�ͱFn�}hz��V,x���<��~�M(H��e�ǃH�L�(��w��צv��AF��	y��Hl�d	�e�~o]�s�ꯟ���5e%�)�0���1�if�/S��W/�
'�]Q���ŀl�fbL�_x��8R\�(��^ES�I|#����G}u�r�b�)`�����zПi�T�>/nB�;�^l�0�k�^�=7�H��쌅����i��/K�@������z�*G_��E��R��*��� �ybV/��#��x@���j�:ʘv������x�?� ���U�5PS�Z�.�q��ㄚ�|
AΖ@T57���d1i{L�{@~�T05���(�^WiI���z��ti��K���7.?��MDY������h�����r��:x@� )^V�7�*���� ���/��O���S�EJf�t���u�V.�41Xܿ�K#����F��wma�O�I� �)��8��=kG�U�ǥ��,H?�Bކ�� Αμ"~�U^�lX�H���P:z��3�`o~E,��u��6�s��p�P�Y��c�:�zw=|�M9O&��6��:����6zV0%,��$�/@B2J�����h�a��.�������������H^��мm���`4�;�O�S:n���Q���@��6������P�ڳ�芿�O�]���Q5�;9�Hi��ҵ�#��}ݒ�<��tNh��7Z/�-�C����sܒ{��$>�h�}䭷�z��v�6Wg��i�sLJ�	�B
��n��ܟ3U�4}f�DY��������.Ӝ�N��N!�
��r7R����5x1��7
,��bs���#�'#\v�U�7q�t�*�Ϸ\NQwdU˷J.�n�6�zK/0�YS�2j�^U�I��z�8���\��*��I�op$2���Kv���Fm2r�ٌ��V�!8J^�������D�M����%-���P��
�ò���o@�$(�Z�F|"���T|,�1�g%\��ᬁIr������#���GY=m���IL���y��"^�^�����/H'��.5�oڹ�ʐv%r��x�i�$|*)�����y#���Wr4�D��K���A��=w�8�kp�zs ���m����7�o難�;vUQ,�h�U��a�M�M�رĵD�-ἔۙո�������h�x����,�a y��U��v���x��!�F^� ^��,�7
S����m�ؖ�']=qL�\E�x/��"+%|�]���Q`�&>�j�����m.��8y����n4 7D�M�e���������r�{H�Kď ݴ�ŭ�;��d�(�5���>)1�o�%	
��v>;HK�����ZI� 0(\Gpۼ�F1!�EG����5gN_bn��83�i����"?��&�.�`�3��'N�6J�����{E���z4��c"����K�M�4�5�)���9ػd���H�A)k����!��r��S�Y1s2]ѝД$�>�v�O���F�{�^��Y�P�D�{�T�@��<��bQW�G��=@,�Z��&E�@�KAwV�eƏ��}!�_�w����\ow����UL����dg�C�%�,��k%A��l0�d1�[�GZX�oÝ+B�4�Ϊ,3-�CVvn�ȴ$s]�<:�(i6�Up��QϛOؼ���orPB��A�nXu$#�z7 ��~X�I�Ѡ��,�8�U�s� ���r=�z�@�]�ԝ-�{R�<�ݷT㍡#
�W9���lq����!@l�)�������tq�ܷ�P�	r��/��)n;Vj$L?�=Z��@ڄ���	Z4��z�������ƗWZF�:�VbN�k^�;�O�/�ً��-��9u�@�ĠV�q<���֒y�m�٦��,����qa�mlӁ4�a1�\D�c�M�
S��>=�D��(~�������,�[`���^Kn�gť�����8+��!�϶�+���/brXg���Q	�F�~:T���	�>N�P�%�
��y�C��Bۓ��RgT��S�Tȳq?!� T�����p�Z�k㼍O���똈 42���w��N��3�^��-��M@�dD+�p"_��I�ۗ,������P�Sl���`�1�.����ᮜ���3Ƈ��}%�o�/\dJ�K�~����Z�&nJj'Ch]��!l�N���/$�]�S4S���%��%���-\��x�;�?	,a�냛�f��hğ�fJZ��Dbj�c� ����z�pn�
�i4�2�y�2��r������7���T��
DU�3x���O�N`�ϽҎ��5�f�ݭ��^{��S
�'B�$3f�bfWD��YmF� z	�֛q�������]&:�������PKq_��v��eFJ�_��X�OB��+��j�f(�`T�:2�J_/��S�k=���*�l