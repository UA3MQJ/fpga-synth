module ModuleTester(clk);





endmodule
