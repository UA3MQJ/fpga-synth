��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>� 0�ʪ�jUаtB��(��K,�!I�&H�;�3�r�<*�0��H:j�aXe�x���
�Â��:�������e� �H�M��q Bq��nwGf��tJ^vQ�Gθ�a0̦�`��Б�0��$��PL8�7��V������{����
�c����x]��2�ݦJ���u�a�3w�J��r�(jJ��TMB��M��m_N�AYv�����������(i��F)c��{{�x��D�Y�#DLD&5��(!4+�^:�F�L��h0e��:Ǐ�*��Uzt�~P�2�׉���<��ư���v���x�&�b RϦe���w�qL��7

	!m��}G�%���B�Y�S>[�H��Y��]HG����G��qF��Y�#=�Y�o��k����|>��d��$����@:�l�$! �<[%�ڜ��]�Ov��Μ�,&pܙ��k"�e��U�y.E8�����JQ��߭R���X't��^��K����k[��<�]����`e�j�f�^�/x����K
���nй���0_�V���c,��Y����Q_\��?u�*Kg5��U�ʦ�CY�q�tlݕA8uX�KB���|x%&�~3&yj��zF"�c�|����ϓ�9d����,��Ah�H����4��m�g6=��O^
�9���M��!a�:ND��d���?��T�5ʒ���3?_��ț�tEW�7+8=�H�������JCW�������a��A���Χ١r3�ns�Ȓ�>$�S����\�4�)�$Vn0a���lM�!����ὔ]ӑ��R�G�����*�.[�"˺���Z��]�uݼ�

���w[��Ԋv(�Ł�z�+���> _��AMͧ�t��Ql�����G��Q��aޒ4��^�4&C-z/�+v�
�U-t%�4��1	T̆�"[����9�8�<�%����D��o�S}�k�A�d�ԧ����V�Z���D��Y�9%�/�W�d1#���P�M�xw��{���w��mxH=9�Y�0T$�m���Dq�#��;�������6�o�
�����d�7Bd��b�1y���9�5�B�&v���πf�V~����s��s6s����W)��9�4S��F�:q���@Eim�Y(ر#���EB� �<�y�l:�����t\�u�K� �{��,�Nh����_h%G2�@�ܡ����%Wy~>��%GbAgIUx���W��7dwR���Bx�U�w��$��@����6��c�*�v�4����-m�~�bl�Ǜx)9_��Y�窽��������T�^v�S��(�	!xӎ>;Q0ʬ�	,k��ң�n^w%��ԭ�*�����ԑ�rbJO�Dq;�YmMx�6˩@��;���D3�{����T��d��C%�BA;�������O����2m���t�h���Oӵ��M^Ĉt�W[�,m�+~P�������cQ,���͉�CwR�$ְ�B��֘"�NP����Z���wǮ���z�.�%���Y'B�up&�� Bb} �(�Q�L$~DeS�ǲ(TtF>��L�24��49n�������B�JJKA��%�{���Gݹo�뇤�X�����E�c�j(�ۅ��Ѝ3=��Y�Ew_&'Ci��/�I�V�} sG%�:�a�L]w,��s�V�wӳ0��r�p�(N��2g$A.^��{^�+�!�?��{���1z}9�E:���=v�F��L������V��֫�M��	��<TWO��)��.�k{F��d�Y	(aO������n��\m�_LF�p�F��D-�zĿ"P/������5�B��ל8��-����qU���?�����_g���4�6WV�p��N��ݢ_�l�F;h�л4.\��=��K잱�P%:\!͞8͋�X�}�Q���;��;b��%�s���4Y��e�(�]Hz�`����_�<D�/�6Xl�b�KW��,<j���A�\�J�mkt�`�ޔ$�ݘ
�D����S��2��4���,f�e�Ԯ�k��O���_�����|�Ӵ�~GU�x�UB�~�v�p��O��z����y����y��cH��^�=$�GY}-���KI�i�t"n��V�B!���']����چ�#6�Ά,6ㅁ�V|�Ȣ+��~�yZJ��6�@����7?? ��\�ꨬ��R��ܔ���3�c�&���_5�Irɜ`Xx���ĸ�&�fd9[ptm�!E��N��ca��M)��>d估��Ҡ���y9O�(�쩳?��Stno��D�$HSq�RC_E,��/O�'�[@ۨ�O߼6�b��\��?��`[��I��a`[���c�y����Ē����h��%H�_��^��?&K껑	�:��K�M�}1ώ��%h�W��E�#P��Pֹ^��>8�-�K��������6���)4�C���&��<��������Z����4��Ȅ�/�h���Q�#q��*�U�sxK�CCR��>1�%����0���r�
�`�#b�`�}�_�0�R?J�u���]tBA���n��38&>)�:D�Je��繷|���"��	��b�Ө�W�L�|��]�z/�Hg`3T����Ħ�p��h5Z�z�f�9�5T�c�w��ώ�R�0�����j� P���'��{�=��c �)Var?o�耊���g�c�W:vIS:6޼s����3���|P�4U������Jo�!.�o�챩��~�{,!3V�Yzy\o-�׻E��������9-�^�I�o��!�4ü��W��ު�0��Ï@�A���D7D��ow�m4�.W�]"�J	�YH<AP��+���.����$l!4��/�������'9�Zk���8�w��DcQ����a4g^2K[s�_�� S4����UZ�Fv���:���A�Um�я�2���G�)|����7>BO�ɾ7/�Tqw�E�{�I���8"�����z>T(H�/�KG��IJ�C��I��a���qd��{��R�\�j�7�q���k8z=�\.�[K�%����_�HU`k�gu�uIc;{,��*��ۿ�.z;<T�����S��K�����a:��[����@ށJ��A^������q�}�	L������*����7�\�=�fsdM��W�9�JF�wm��n�W��;�Ŧ��W.B�"��t���qdSͲ'��(_��T�~ݼ��R3������C�L}V�����ψ��!6HXl#!ڊ�s̈́JSo�Pȥ<��۠�� DP��E�sZ�#Wb��20��g�=֙4dĥ�����x�.ە�"a��12\�t4�:='5���J������h�7���