��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�qޛ9ܷ�$��{��>H�����.�o�9�5��U���S�FhuA�f��GZL����I�yq��V��X��U������~�A2�z4a��0�L�S}˃��FG*2lH�M�_�w���nRl�'����!8	��_�/鯹��h'ι�����H�'���g�fXR�O�v%iBFG��5k�3��2�����2��B�M�3`𒍧� ��G+N���$2�%f�w���P�����(8&��"�
�d�3�!fu\΢��h��5Y|:r�2���|���Aoo�X��.4�-���L�䌈펺X�z׳a��h
��{���8k�֥�g�D^��OW�:�d��P�*%����hM��~㑍��6��G)�.��
�Jx�7Q����s0�-\d9�;bY������-L�ǘ��,Qv��F�L�E�&,0K^U0@u6�}����:+$��6<��C�VlRik��wQ�z�T]�,�(ݸ���&�������^	RG�E`�A �n0�r�"��
A�&��vĵ�o&ps�����xR�Q^F�8HR�E~����]����"���`���I��|�����W�RG�c�v���X�O�2��AP,e�-�#��oW��}�,U�"��Rٍn�~(���0#���7O��&����9�^�hʭu�t]��)�O�
6S]k2�b�_���o��LZ��v��+�W%��� 6�8�y*썎�'��Q��ɤK���`Qۚ^`�
&��v�D|��|�$�in�O���$�iD{Vg�(f_��{!�L܎��\PnT7���`l��+z}��zlؤ�E��}�ze�r�/J�W�=P��U�ԐÀ�?2z�ڭc� -9&v��U�c�Ŝ\ek��g��0t,-��.�=��s �u �G��������Ka�H����@'A]>����$\;Ydv���1��hơ��ޱ�6���a�uFN��x[�zy�)$��s���@P�D��#($wn_&$����nj�f6"/;%�?i>�$|���������I%��2����O[=^�R�T�n*�k��F��Υ�8:��L;��s�A�>@T 4��G���y���5|1pW�M�J���y��@�c�E~B|�.��E3i����F��b��z�i/V[{�~�0~���*Z~��B2������Z��a�ܓw��vG��z���u�������*���NJ�Q�ǵ��M��̑���'����f#Z��D����\.E�ƽ�<C�G��4u��G;�[ip�K`���&�Q���r����f�Ap^c++3zEb�mmo?��7H١GG'f��7t�m��X��Ӑ���Lxss�K|s8�W���O(a3����������L�V��zNJ^����>	gt�ǗX
��DHtykH���+u>�;��!�� ��G��U�ܽD���y���q�D���ɦ�L�g~1թ&�q*�s�:p��6����~��r�/��f\�a�UY볅4�T3LkTV���B��r]�����kr(i��+䯫��A��y ���
��!Kf��ȧ�#��A�J�U�j�i||@G�Z̢���y�/��D�ZE4�V|$ө�h�����Sx��r$U�nk���^ݙ�,k���.��nWy_��}=i��J{?�����Մx�o~V�w3m`�y+���v`�CPK����j\Eo֪�V��B�Xޝ�x@���"b�j�i4���ë�6t8�0���p��N$��Kt�h&Zw�f뷊�����`�����\
���qܲ8O�Ȼe�0��Qor�W��M@ִeǣ�]�$�z'rL2Te}��/ʘ7n�N��6PC�Fx^�I�3����Ug�i�r�o�{a���[u�	����]6��c� �����=N�}�7J6�>�D�9b����d߰ �����_ �&ٷ꨻"a8��v/Y�rk��u÷�ՠÌ�%&~2CF�m��z~��^�z�9x��,W$_�N7����c���z���L~��wSO��9��[5!���Y�^���a�Z}������)��x�ӈ��Zo�2��E��Iӂ}���ٲ���)�R^<�@|��3_WՄg�Wl����g���c{BҼ?�["����j�ۙD�b�����R������429�@<^������vS�ysoi1��kP|L�p��*��B�)X?�)$���>
��4AI�l�Յ�FjV�Mcp�&�k�h���i�#��DA�˔�|��J��9�7*���_�h�{zz@k�O3��.�n��V7�l��t �(or8����4!��@V���ܓC�wt;�p�nx�9R�7mg�3@4Hm	m�!~�7h�B�X��.b�Fp`��0<� h�Ci�A��r@p�5�U�Fl���2��r������;����!�QBa衑*ݮKƕ����*ꏨf!�����"| ęY��o:��u�� [�8�V2>/o�6�^e2h1�4;�oeI�ڭz�c�`h�A qv�(����:J>�Ʊt4w�9.Y�4>�u�Q�J4c���c�|)=~��H��Jnd������Tc��������5���%*xvآ�����l��Et�l��iQLd&�#�Q�H�L���WUc�-vGP1��I�Ӭ�Uk����YJfl>Vy�.�M=fs���?n���k��X���}�3�^4�E�[T�2�9�VG��6t�h3���jʧvN����z�oK��| �� �U�]�u�Ճ�y�F�~�Q��2s(Xy_WwE�m+?��Y���d��<�x*^U��:`����ڏ�H("�bŭ Iv>c��2):�cd`ԯoZL���Ĝ�%e�=�wi�{�[g�ғt����T��~n� o��PFaHĿ�y=�0Ó����\�w%%sQ(��sr���Z�����r&i��ؔ]ѻ���V!�����wK��' %�Q�S��:�'����g�E�|I:����z���� �A#�W�I�#G��^��Ƥ�T<������d���v��z�,6�ix����� 
�a�h
�#�g�E�xz�*㕳��m�Z,��.hUI\��B���422�NԷ����}�!��Gb��h)a�A�p�ƃ؆��numqJ�]$J��;4����p��k$�H��H��I��`�*���}hl~�(�����壱��sf�"�T��I�f��l@��B����xmȚ��&��J���.aـ�7�v+af�x�s<�<W��>�܎6r=�>a?0.O�}�+:��AIX���%^���1�s$P�&D(���$���?��W��#Y��l���`�d�v�8b��Cd*�>z.~hQ���*��X-