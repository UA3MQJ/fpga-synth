��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��l_����b�-V�m��mZ|�)}���j5*�q\c�0~���dwg[�$���ט���N��Nϋ���Ⱦ�[���|�������������Ҟ��(H!����qr�2*t&�![H��Eh8��E�QЎ�D�.�(­3���b���Z����L2X���x覑|�c)in����=���|���V��`wt�1�.�-K���,~/�S��3Y�2�QvC�k�Go��#���#�L��������-֒�Vд�NN���!�9x2����?�k�X����]gM_�h�7H.QWQ��ߥT���g���
��`�	V�}�9'����|}�յ�CoXz1]��T�����p�<�K��4�;��9.�&ǣ����q2�_�������oB��1�3(�#Pu*$KK����r+����Sy��jdqڳj]���j��㏎�Ƞ@�)g���^����ZӨwr�yBp��˚y r���.9��j� #��'���U&���x7C��߲{��&Y��s�ew�X$���	i��)���<\ʦ�۴�]z'�H9�e���J�*�v��,��8j��s<l�)�xf=���9o�wɔ(���� ���L�2�&�}��aW�cl�w�_��cOD�|9&�/�5z%h�}54E;d���Md�x65M\�r.�gk���H��+���B���L�/���4'Zt�t���I?Vy6i1_]���-��6�M�Al�W��tr�h�^t<�-l�E���C�*��s��������@�[_,U4���b�.�=E�q�5�<��qv��Ή�MP������`
0;jz�N�>����wMK(ȸ'�T��D��s	~<�#)��3�cm#AN(`�}
A��˂ �=5{�?�O6|{�n��ro,ƓP[ߧ�*����]���$�@��W��8ߠ���1����9h�c
S�;Q�a]Wh�/ш�����\jD^��{|t���(/ �y�����w9�]>�2N%n�e�~�/�r�nCY�U�}���);2�Ǵ"����7��6u��G��-Z�f�6Jͽ�ޒgc+����t (��8.
�[�~�Zڠ�)�evq���ZLZ{�c�c���0Z,K���Dg�6��^g��Q~�ܥ� ��|����A�v�&+,��e�ܓ�l�P�A��3�-����X��[M�V�9)��K�#*��@�6EG�K𡘸�
ƾ?�]�suS�A��3`����9I�c
:r����QV��N�lB���f��S\�tP}&�7���+ /�\\cqo�0e<l�zJG&P�U�\;ƁrG�_o�^�
Z�p�A�s���U{���r�c(�G<��_KY��H##�Ѷ�'�֞�������#�it�������D��8�p������=��P�l�78��W���Ý	�ڸ����md[����w�!5��IerE	�u�<�~.�@��dBPC�[�D���[��c��y�(�9�?�:,f<%��*���� �R�SH�QT�T��m%������%��.רs
�O�&Ջo}}0DzB@D��Gcp�(.`���`U��.pIc���l�w*[Hǟ\5��}Q&2?�{Yg�V����ZW����.����T�������ȣE�i�?�X���D�/,�;M�$��.r$�y~�D����#��ުx�W�3��R3�*F��o��)���[A��z��o���f�£)��b�rϝ�oB�0ޥ�����,$�!��Nw����f���2{JR��P3��۪�����nƆG$�Gc2&���l����thF5�X�U�p~�#7�����<i?3��?�p����'ږw�@犕/��ǹ+4��o��6�J)�(uF	������c��q�f�*ۍ�J�,�x� ��7~6c�2
�Ra�ф�ǁaZ����.*/�)ǯFWH��ٔ�u����aPTO!Wt�4{(11�b�i��D}�"��%��G�[�͞���q\>�1����i6�M�|�׬@���^[]ҵ6{�`��{��̩�2�$��&�8_)��{���;�Ե�#Q��q�s,��8b劑�@��'���b��ĥ7��#���4��`��)��_/=B�Ա����N�6�o�WO�@_�N]d���x���0��L�Mߠ^z�pf���۩B�:��:۹`L���*�du�ѩ$�i� �`�`��s=D*�ii�}�ll�"D�D�U��9[];P_�"+���u�Cq�`#�~	�o �X���C~��ү��m0�����XJ�d�=˱S$��ȅ�ũ��lA�k�u,aIl��_���A�������`��N� q��=�����e4v�����gx�-�� ��E���S���1�#a���ܮ�Q�N)��yBR��x�/<v�i�!� P��OɆ���ґA�ɸcف�8J���\�gC��>��������t�}�,�E�ݒZa�F�F(��\a}h:c�����W"gL��M�Q!=�,o��o�e�&]�C.��J7Ղ���0�JaR�^��/�8�:��� �ȩЦ Cm��Ĺ�R��k�W��t�B�b��E�I>�%�mW�R�)s�������Cs5P��q9��*�|8�u�-[:���y��|_������ ���15s�V K���Ff�<�٘�cG<�|[Ls�糦h��u8�y�:�i�G.:�daPY,����#9yvթ�A.�ش�
��IF��Z��7�7<`�����Z�E�����D�"Z����� �|���<�_"��M���֚롆!+�וm
l���*R�����`�38�04��z�j�n�]e��1z�:�8�ϫ2������1������v�@ʱ*�:���Y�l^�6��d�Wh+�}�jZ
.I<�.P6M��G&i��4�m��@Ƹ��S>u��ՙ������}6W�Q�i��������誽�9�$�$vuӳ{3�<���9� U� �W�U���&6�`缎�I׼H*@s�j؊��K�"-��r��
�0�7�2��yǃ2ڼ\Gc���Q�.��T0,�+^�" \���A^�9�;yO������zz�D�7���~��\������n��4�
_HaI��ߢ����l�G�--�O������{g�X�9���j�>�.��m$�"�;Ӗ��O.s��@��������<+���n_<7V�DQ�H�]���&��L5�|�%bW���H�X��l�CmN�aT,p������������-g8��_���)��6�M��ey���=�-����y�Ks�5��22�:�U+�{��b���!�Q�8��"9�AX/n71��=XR��\�#��Ϯ�Q�rG(ZnK5��xo�m)5���k����$rk��nf�����ş)��G�=� wX��|D������F����?�"9b�5F�H�<�B�0o��,]����+���n�ȿ]����K�����X����&!�'��6��?�������'i"�&ؙ�{7�6jj��r��l�^��xC`GFX$�m(i�\`D%���|f�
/W�D�H�:�E����
l�"yS�>K�ؾE�*�Ֆ�;Wl���i�:w?-���g/ڢ{�g�7V�)�5��K���M]��,�T��2�r��U��thX�MC�&��a�k��W��{��Q�@��`l���<-����#ѱZ��(�\?ҧ}�Iq�v�(�������L��)C�S��Lg�������.��!�D���G���/�A1�����+�K"r>ݤ�v%NQ9�D�Es�S�,6l�,褉"7B���b�'��3���4���.:N�!8���R}��|XT(n�K;���t���U��l�?�^<U�5�� l!�ON���bbƦ�z� Yi��݉]��ο�6��S������n���|��!``��w3k��)��~�O$O�K�O��8�*�����6/�h ��,ޏٸ����x\�N�לhr���m^�A�A��	���w��;�KC��Jb�6��S���'r�����@Vg��]
��Kk3��)Un;�%�+�x�ݵ�e�>�=���T��Ot�F���q��f_��Xv�B��87�Yi���DX�9����
��C-�_N�9%�r#�hG-�Nye*0��Ƽ_L�nҁ���?�,E,C�7G|`��*�����e)nX��մk��9��Hק��N�0EpP��y>����].�K6u%�pѡ+���޴�P�r#�^����4%����̓uk��'P|��JF��-��[}��@:��|QI`�kL.�+Y�r��7�$��+	\߲U:G���Vh�6�Ң:��� �\7�q`��Mm�/.f�o�r�Q�Hw:?�m����á��B�\�1���	���`��JWv��~F�,�X��^bQ�R5��]GA塐 �U�*�������9�W��k��VSM���z
[f��<�U�^&�i