��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4���"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!����� �@���4��8
Km�'��W�t��㳥=�,�Q�{�J,�V�(-�&y�����+�I*-h�����'}��"9�#y��t��J�H�.3]T?ֵ��#�C�c��ҧU�d\��2/L�5�w�����?������Cę�,��qN��I�b����7�g�#ɧ�-�u���l]d���*�|��*����~TuD��ܕ^��V�.?0_�#5�8��^��j��O0�HQ��oo��U遇Wزk(�-W̓���>`5	��F	���ϵ���}��A�(R�I�Aa�¥������e�'U7ث�I�ĉ��S�v�^-hTM�C�i�bSk������g��p.�R���T�Ogo������ퟪ4\�;p�񾲞
�9
�B^k�M�X��`R>�dW�-v6P?B&�]QTT�ve1��'�7��H��W-��b5=e�)�P�ky�mlL�7��6�8I�� �`>@��Y}�Ŵ��ׂ1�+Ǹr��Yf͕���
��)�2?0��́�&4T��u4V?ŋSNq�^J��r,�| (!%���^'����
9u��J
�&Zm��%�eD���E_���v���w8o0s �����>Z���X %���Ȝݸ_�97��,��Q>��Hr|f�v�� �šM��'�Ԑ*v��>�Os�\���=u�p���dbXX;��l����T�����g���C�@�9VR�MӔ�ZA~?���7ږ��N�E��Fry��`۱W}�*�7I�+[W_kO��z��?�јwr�%tl�m�lx��M�%&:+ͩδ$�`�Z�2|m�ثvHS�w�������>�P��u�|��Y��"�q�*��^!���d��	���v�K A��F�����w��	vG8�t�@]Z��q%�����lʖ��݃�b�[�_���r⮿��YJT��
H_k�ұ쾫85��[�4����4ô������pU���*��_L���d�C�(@���`a}��+�	q����:��n|By���>�N�:Wd�^P�:n?"��5M|����T����'�NV�5������*uya<��J\��9�o��<D8����m���`×,#Gy���u>w3P��&�ۅ�We��t�%��c~���j����6>�H��Fo��G�.��y��7]�jX���U>�ŝX�l�ԗx�<��2���h�kU>o��o�1�~f$ajT�"Ҙ��F�)�!��7��G�rK���s�}Cc���U!��G��.�@(M��b�+�/�A�x���؟D,���ɿq{����-��p�q�%x�9��X��9S����ix���S�M�+�Δ��!Q�L�B58l��|���FKzv� �,�d�tQ���E
����1�K����*
2�]�h�Wzfp39�-�(^�o���ו���.��J�)�,�{6ٵ}q�{˥G�;;����4��9^K��%�K�62��aa &��,U�R���!���t)�$��h��t��HQ�Q�zOg�����g�k�y���m��ڇ�W[V�S�J��U�F�c�|�=���gt{&�[�֨mL�!�����~E}5�����Ø"�V�	�j�d���|�'�\0
1x#7ͯ�r�Z��|Ot�&���M4���J�Ɇ��~!5�2;�QW �`���Ԅo�����DU07/s���j��Յ�Vt�
������|���K��<Ca^k�ǃ�
x��A�@�9�T�An��*��\���U|��+ñ��7M�{{�l)y���	��[�j�e������K�VJ1������:�@�x.D��,䮢�'���w�@���$cu=��l��٩�V�fh�}J�1�鳊�I��+�@["��4��:��a8��y�Q9,�,��5���`}�N�UwU�|�>�`�6�E49̖���A�2㟬5rg�OX�������a�:I���(�Ы]��!��iH�MpJ���u�|-�Σv~5հ�6A�H>:��d��W�&��<%��s_}�h���H��Eԏ���D;���s�O73~�AG���D�瑀1K�t#׾��Z6�Q+݌	�4����.'�����pv���yA�����K1%�O��.������"�;:����q�d�7��*>�Y�VѨ,)l��&u���P'�'v�
��P�A6�;�>%kW��n�)��M�WiF�\%FrT�ot��_�c�I��*T�&��G˘9�N���U"H��؃1c�x���������,ƹc�V�M1�^����_�^� na��1ѳ�픍qK�J���O��n!�>��&_����4k�춐%,��D�3t��j~B����5&B�+$�P��?7�����A�:]����=���J��g�ـ C���RlTj�92�L��[N 3�T=?���5��ªpE��+\�������(�'�mx`!�"hY��.��B3�2{���� �,wX<g�X�(����a �uKO b���U�������x^��pu��L�3��kW��W�|u�4��g �@<���6���Ƕ^��\�V�@�i��>îW�pIڄ�g�6�箤Z�)+y6h�Dlh��Z� �$5� ����<4�T�!`�� '>�J������>��^_��z��;%�̙�[B���ǈ!��O�>"�U{�K��d1��̢��EC%I��Q�������R�_�I#�Mt�CS�^S�Db�b���t���X�� �RV�z�y2 WD�ΛY�/�?>'�]�IU����)+���S�R.D�X��>���Y�˴R��V�ƨ�5ݘ�G���qV�Ē�I�c=���: 0,�����>��%R3m�xל�꧹s������s=Lm��x�{�pM�%q�c��vb��x��������`�P2P�p}�QK�S`
�֚1HЅ���C��!�r�y�,�.[�l��懼��QQ/x�8�9�/�&��~c���#�6��,�+��GA�+�׀HdVYC����bI*`�ˉM���d�n�Uv�
���5 ��i��d����S�� &m�:p7(�΂�N�h> ��-ӝ�4��nU�l��eAZi���B�;f��9��^ R�>���g�w��uO���ؒ\���7�D���ǻ����8aJ�c�V2�y��Wr�8��<փ�sq��U^i��|�4@%l9�w�c�5U�T��C��	��)N�S�|�U�z����sD��v���M��6^��Lɫ�S�*�����\LK��K��֎���4	YY�5x3�G/ժN^�IS�/�Ц+�4�x����m`n�d�j�MQ�~�8f����Iٚ~�2�O�,�kl��}n�/a��m-q`��~?�k��u+a����M��_�2;�����2>C�{@+�T�J��~���΄غ?�	|�M��xy�,�8��)�4���%�_���5X9��qY���VF�o���EU�뎆�p�eoQiQ�%���]cGb"$�z���v�	�4�l<�|�(��why��e�"}�Ƕ;f��⳩#]/�M���j�A�1z�i�[=��;�X8z�d��0>�f��p]@�y-��mR��o��t�GJO?gJ�k<��0:�������� �%��~��}��m�}#?�S3�v����I~ a���D��Iƿ���X�ʡ;D)�8�:kF�x�q�;��p�=w���0Z��WV�O7�	^T�'� N	&퍐pQ��*���,�S�fz��TKÝ���u~�3��h���A��wh���Q���2�A����Z�1d���9�Z F&J�@��q�^"����.�;��ۙ��30�>������7=�zs
��\x����c�9rj����GK�	k(lnchq�u}�u�q-e��?:턌M���Y[�h�'�rvjQ��U���`}�}�,�Js�p�P��eh?���:7<��ofDU���x�����Y��4%�ݩ+ZF�DL^��3���w6����{K�A�y��R��A�z�%�ݪhe�}�9lY|Ŕ�I6���"��Q�%�d�wߢ�F�J�}��w�.�r��)8�Zy�I�ήMsS,5�]���3ƽ�I�&ԡ@��0p[� ?(3b�NG��3�#9���9f�$�X�)��z��ʅ�������Â	���*;�5�ԁ��E5�Ɯ͸�����6ݨv��c�n���
����p���&O��E�ױF�f���"#6?�R-�AhA� ��s,`����)!V��c��9#�u1"���,��?i	S��ptWx��%i�p	�2�6L������%Ti��'n1�A�;pvcWGɅEH$�<h�����娇]�	�8yo��S_��C�GF�(��-�h�I�:��I=�V�'�<Q�+��sCμ�9(랤�~H#K��Qd��H{kS�y��Ra�,F.����Ħ�~z�V5�'=��H\�[x��Q1ï��:Sa7eړ�:��A�x�MGd%��t�6�]Tŉ�up�����J���=DJ>�5�lZ�lq6hT�F�J��������$�oQ�	�2�j�>�Zè���i�7ֆW�j��8 k���v߹�T����/y�'���ӏ{���Kln����t��"4U��}	���$^۠|f(�������G��ZtU:el�����u 	3��j�\9��b�b����X.�Y/���1��M����1@��)���o#�2عB[�ٳ|�+���Н�YĻ�71�����]u8���%�b&��%Qc�[(�W���[z�x^:�tƵ���� C2@3����kt��	��L��l�`
�J�'�i�d���d�sY�d��&*>�J��o��DP6��v��7�}܌���՜&e�k�¹k��	M��Qa<���� "`��@�-A'w{i���PݙY����hf��g����d�A�`F���3����`<�/l�dt��LvX���Y�b[�++��_�S�1ԝU����z*bbם�a�5�˴ރ�z�(mLa�D_�k-/J{�%��_�N�a�&��{+��N�:�o4��[��Xב��8�+��t�B21����2T;粒������d�!Bڊ����5n��=)�`J'�(�FkLf���4�����̔��D�ŐH���ܠK{j=B��"I����LqË$9�mA�]�����J^����r���F+���4!�O���}D�]�vnJ��/:rJ!x���b�����_T�U��Ya8�2�/�A{!��h�$������o�cʮܽ?����;��a+o:hdYӌB�.�p$�S^7X���8Ƿ��+�ڒ]������������lB�IA��Z�-6�J�':��l�X��ʨ<���(�	��K���]����iҶ��~�t�;�
�=-T�V�oM�?��X:{ꉞzå�v% ��@��mzR�~���im+��I5P^�U�Z>��vB��)Y/t�_�? �S��	<͡�AxH�����K�@���a��DuY�1��{��\`~���|�/>R�JaD�i8�6��p��	eR��5>�����7�k�pE,��5�h�.�@�uH4�n���^Cli;T�X\�69�������5<K��;�(��L5��l��N�,b�p=�5auX#�.�R���&���V�3�#T��cB�h�d�É�(��(�qے�� ��X���t����c��Sl�cq��)K�����ޒ.fz_���jFIj�E��37�сV�!Y�S>�s3�pN"˙����v6�b�m<�������]U���ǁ8 �fF�n���mk\�>��*�*..�P�P"�nl��k��o���������+Xvy�
{#�%��ػ�\o
��M�%"~�RuJ^zX�"F�o��,��R��c3o���\H�ꮙ7�Z�@�:�?»e� ��>8a0������BC�/FZ�o��ôB5�}i^ /�
�e�`��nP��2�֨xy1����<%��2�9��:�Q�$��2MZ2��W���3���1�g7�E^����o��}bG�m�g���<�;�{L��A�X�{Y�d�1�dslG�F��B����t/fi fʹ����K�q1h_��gF��l��,�~��ZhĖ�d���_�euEy�)������R瞒���(
���|>�6���y3��T9C_�`C��7ۄ!��&-�F%[�>-c9��W��I�Mh�4� ��fgK>+$�z���u~�h7?ݖ�E�,�]�H�ڬL0��k����\%g�4���+����S�mؔw�o�5���8�V$G���ܦ�=	U��A���+o���騚��j��Ĕ�� �"o��UJ�$�U��t2�uUY-[㦭_#��BR瞚e��Ĩ�Sg��U��J<ٜ�T
�?��)!�ĸ%��m��l�{�f$��Ȋ�W�ӽo��`����=�[G7N�dyy�Fy�ە��{�>�,!�L\����݇R)�HS��+��6��3����nHG���uȃ��,\���ƏtX�+�t׍Q7N�v�L�ߧ�!�Z��y�!���.�8�%/;H|�i䯩�����pl��(�c���r��KU��Ħ6wK2Xd�*�I��U@kY�ܪOu�W�J�����#Ƣ�.�%�	�6gtMRR����� �a =�y���y���B*�������� /�bcA*俤�;Z����hz�n0��:-�W֌n2S?����~�%-��e��B�
�a6V�S���2a�sg 5�Os��E�\�b�|�(]��'B[��E�&B�_�CW7�L��wl1�:���"
���M�l���mgwC1A)_�<� ƕƽ,�P)P��M���ͣ�|���gd�b�8i�q���G�ş�(�������}BAN9�zu䥢��X\-R�M��"+L��X�<t���dT��M���[��T�v�bov8K�%�A���1e�L�bhω���B7��z����HW�Z4c?��+��u6^�XS���H�|�W��ulєb����G!5u��`�<��:��p�lKV����uO�Ic&�,�#@��e�*�"͔���o ��^�B�����C%�W�,�����S�CI�-8!��d2���E��;�S�Q������c"4��
�)�$~( ���$eO�� �lR�kAq�����Tb�
dەh�o�`�6�\8ݸhm�x�R�l��q�F��*-�Ʈn�Aⴥ���%Q	Bр����}�λ?���*�/�g��gs�˼p���t :B�,;��~�V�mri�{Kqڝ�����N�%�҉�2����<Eΐ�9Ȼ�����.^�����4,5�!>�2��������:�2�2M����:+��K�T�$'1�fm��}*ei���W��Yw<���H�ł�:;xߞw'|�f�Ip6P�."�'}'2��7��qke"����Ҧ�̐,�����m�a�\�z��[~\����YW 1��|���~~�d�ͽ��/�Q��V%N?�#��LY�?�j�	��\��D�@�#��Zp��A� 128�l1�xLj� L,ԓA��SV�b��VwN��|�g��RW���22�|׭�bmڍ�̺"	���M*���U���u������~���+����}�V4���#z"��3�Li�������*��`�h� �������0o�?�lӑD-�>�z� O��4�Q%U�4�Ƌf��Q��HK�M�KP'�i�Md�A\�A)"��j��_j r(�n
1��T0CM'�g���ӣP������Ss
a\�!�X��oPܭ��1ױ��
1`��� ɱ4��a���8�y}t\�UD�8�^J7	��Pr�Q��E,������`b6��Ad�8U�>O�q�<1�ʴO��-c�T� �[���X�q�J�,�š�(4rF��*�B׳Ͽ0�6
�?��mt�ı�b��2MUhi�7�ۘс_�i
'�wT@�`[Ѽy��Wkw��3�nxef�;4A�>]c3�s���2��u��'�E�Ѕ����xۨ��X*��-2&���	~r�w��ݷ�q��FN��\��/O��WA�����
�o!B���-f��OWL��?�2q��Q�s�K�j4J�@�>�p^�Y%�Yɇ�t@y����E�Zl�R[�_��P��4���h>a�l�sE�x�t�[��B���)SŅ1��!@� �QzEڋy���"�����ʮ�-�Ͷ��2l<�unI8xhW���G��Ò>3-��^	H�����������D.�r6ڟС��NwoM��ޙQH |>�K��4��v<�ٵ�{z�gF���w=#��$�@�����<W����vQ@A�4)��W:�E���qAXBaf޻>���[�^�D�X�t�Ej{�2�>,�x�`Nq��A�Bv|�.$�=��$?egƦȠ��.	e��˸ŉ��n�'cQ�}9���mn�J���Su��{8�D�HF*�yXS"�Uϣ�+2FQCA�R[��Oznȫ�)��p�{?#�]ǲz��{l�t]Ӎ@�=�D%�Q���b��� ���v�pf�Fo<{�jU	�>�a�x:Ȯ��6ƭ��~����<{K��;�O&N2����$������]�C)Dj���5���(sG5lZuvo�rih���*/@-��V�.���lg�x��q��.n����{@��I���@Q
�4TZ�)Ǩ�{��F�����\�l����P���T�ZM]�[��Yۑ:Mu�l�=(�_)Z�p�/�i3lR�$3<��S+Bi@�n*��e�7�N����so�D/ ����u��;}L���Í�����D���I�*ڦe�>,�2�tJ������-͡�BMو�����+�9��ZV�+�̇��u�eH�m�{�Fvk��:ăn�J��I@*�`�O;OV����c�a%�ɭS���r����h�$L�;/NI�(V����K�) ���H��x{H+P�?[v����&L�}r��A��ǫ��gw��sL�@��B���Pl�&n�f@��j��Y�DJ�C�&:��+}�`g�D� ?.I�5���&y���=�����9!�p¸%h�X���ڢ��H�4r��T)�s40ԓ�Y�[�( 4��p"#zK��+��ơ���J����Ne�a�?:��)�Y֧�� �r�cj��,Y����~��k��D�po��wX�/�����W�Ӗ51'm˘��ȥ����Æ���y�fͽ5�5n��̀,6}=��@�^S�m���SE6�#�DcJ������Nd�>�m
$c���2/�y2o�L�3}N|�� ���Ԛ�-M[���C��� #*�JxN���'eΌ�4=郎$�?�
�j�ƽ/�j��(5��W��y��噊繁{,��8�������VqUT��oFK�Sz����t�ݧ6�	2�؀�	\��N2m��/���.�ɽŕt��m0X�Xʹ�۰I�ZC`�������5�lh~�7��S+ޮ�X�:䃉׉䘜�޿�vΟ��u�M>�I�
[}0ah&�hVp����
�?baz?�r�ڍ���c��xy�SK	V�X842ֺ�c��~:�Dt�FyDm9�8r�p`"k�)���)�3 ̲�Im���h�Y�v�J��}u$'�4a�t9���c϶����;�s��2E6�C�F�}��k��|����nw�UX���{t=49fRSƚc�Q�Tp�B6Ű� 3�Anx�n�R�ߦ7����G�Ob�1d�IHd����%刺$�do�q?�z7b'�����jŒ��%	���"ڃUWµ#�.s{r�:f���|ߨ��#��� $��n�Ӿ	��G�D�k�z��U%�&��[
��r򴒀�Y&Æ��k�җ�~�>�������\<.M?�]O�=�L�G�;g�=V��h{��3�<�ݯ�A��8������`�,�M,����z�p�]��H}Ϳ�9�8�z�K�������x��h/�UDl	/��xϞ�q0��QT��;��ch$w5�I�B%�%��(�jXe�q�{�˹������D!�	95����5=)b�f��{��H�1�ete�v�vZ7��4%X��)gG����e����"Нl��e��㊊�6O(FR�Y$���=� �:wNF�Pi��NA9�X�s�A�M��o�{p�Q������1��Z��fJ�Fm㑼��v�[%��M�[��&А�E�L�����.q*�d-
�g\^	�!׊�|���T~��v�e&!l$<�@Hʽ�/��8ӥK��۵?@���U<�"�\q;E��Yn��p}�,[�6o��U���L�.���}�iɦ�S��or�Nlq������b�{`��ʟQ�ɯB偭��h�� >���{J&U�e��˖����Pb�dn�e�]lF�CRu.��aо�<Y��%��0s����7���g5�2���7�����pU�6������r]�4<|=���jns9Py�n�?��S����_���Ft�(��Ϋ���SH���};[��{��%�I��d�Z��mu��3-i�j�w�},���CݧX��	0����O�(o]�X�Id�| �n;�Z%��l�CK3��X�NӦXnЁ������B3�ޓx|׋���b+�X�C8�[��V�ǳ�cz�]�o�і�8��V�ɗ��z�*�@�M�{���2���&s��4�n���b�H֎��w�M=J������,:K����5��6�R{�Nl��9�#���h��,~�[U���c1s��w!�߬R1� �pB�'tڢ�;���?���#�n����e����=�$�O��r����Y�φ���WB!�NY��S����th��>����$��Lq|e�hO�=N�Q4^�w<w&�C�K�~BC��ҏјq�P�܌�1�X�>/d��)�o�&�/h��aAҰ���	U�X	����g��l����1K�4O�L�%���:���??QA3���E 2���]�������|6��΢��Ю�qf��{�%b!�K_��4'e{���\^&�2�������Fv�����ŮB�z9��<|�PhL�B��o>օ���Լ�:���=W�&Y_� �"�z���Ӳ�F�=���i��v:�^�9�"DU�p;z1�HZ&�㈢m³��
������
,�`h.���bp��V+u\1�@�δ�g����Nq�%8��ҷ�.Fۦ��[?��z4�E��@e'2;�M/Ѫ0J����1�=�}������x�p�{�|a�U����Ϥ�CwAB���8ps�G��b}��.G\9��h�4�X����u��H�R�ߣc����@��X؜���]�|�x�@���-��	����aYoe��Q��r|;M����hK�ۙ�j��ˇ���7�ض;���fw��*��> ��E��F]�C�+�A\x��g=5�ʚ׀�/�tʕn��3_w�zQB�i�U�cv!�\?!͂�U�jӽSmC�T/�e�,1[���X�5���heJ�i��/�QB�Seg�H���[,L�)06Wk}Z��ȫ?������:dz�:�^�}�x�ܧ�Y���e�oJ�& ��P���|�����SF�1���#��NI#���|U�΄���_rByG��@�MC�$d��4/��u�p��W�~�w�fF	x�zL�B��#-QOY�g�.����G��p��]�F��F�J!
b.�e����ݐ�hn�7Эzc���z��iy�L7,����2����q�W g�Q���$f��G�.(a���~�����.hVZN�<�NH�/&֐�G��r`�$�Ͷ��:���*s��YĘgr�ʬ��������A`ą��
���,r� �ؤ��D�3���	a�~�!�qM3����b������[=ރ�4d�wb2b�GR�,�
�}���!o�ҕ�o�vO���~O��XU!���X���rXg�g����S�����eۼb��j,�?��$��6��3Q=���I��^��(�rp�,A�C�D(���zE�����Q ,|4ϝmŪw풚%$�2V+
:q ��ĩ
�C��O���}+O�>�)
��8�9�z��|7o����M�������w��l�V�sMc���.�ؚITʌ�G�GC��Vm1���:ډa�����O�
>r!3���=cV��1��j��fJ����rL��w��{(i+����G���s�
���%K�a�]zְ�ʅ�z?e��zlP1�1د$����Hì6a8�r����l�u�6�U)KAkVA�!Ä?�j��4�c����!zG	�S����I�����k��`̩�oE��3pk�5i���GUe�@sU����)����ޤ��b ��WM2�JBn���<�{��Gx)g�(���tZ`[�����>.�u3ʖ*T^GeM{^�e�7m$��QX��,w� �{S	�.x.�x�������7��ɤA��^�XY��c�� �k] L&��R�6�7,�����P��pR���g�n��ҡ��r_�mڀ�B�ʋ�����0��hfT�"<N[��sM��ICg-��ջ��V��\�;D�eyV����J�|���MrS�aEg6���cbY�Zv��tOM�j^����,:����]|��c>lD��$J������b��(�J|�w���jDrJ�U,C^o�z��L�����ED:��U�ī�����u?4�`Ց`��եY�� ?�հ��\�I�y��x-�	�0`;9�/��V_O�ǷA7'#?#!�r��xEN7̀5�=��D�%?���$b)s�FZ$�U$	�^%�5�g����uf�K�b� U|���WW�+�'�JT��mn�}����Oɇ�߀e
�^�3f�ˆ�K>�|v{�6�]䣎7wn(^!�ZV=��y�
���U��>(Ui(��ڥJbv�jW/rJ��]X���	w:��;�!׀�0��3p�y�)���'�
R��6��/���?�-N���10a
^���B������a�P�طd��<ߔM�
R�r-�F������b&c��	���֜�s����+�_̺�u���
���G��3��1W4X㗡��b9�F:�+�C4��d�j�I�wC"��Zu;Z�f�|�'��*��o��t�X���i5�C��{uO{�
�+v�b���i^ B-�ڈ9�K��V0`:�i(�;��m2YP�>����h)�k��O*�Ϛl.�Fjד,��E�V��?u�C�.Ţ]�V����o�2�8�K�é0f�u-��8�y�x���~ �T��ok+�x!(w�J���<z�o�Y��,`�cKVݾ�E�i�=��#;�q��
����5rG^c�'Qs\���/�3��ڪ���P������f�U.oB����>L���q��ЊzbI�[�f��u�('eW~?�(�Z�����~��5N����Ąx��-��y��w����O|��W���� �q�"ψ�@���ǡO�6u�5?�m�L�tN�~�y[��2�``U�&|�NIY��z� �ܝ��r�.`� R�y�u�q$X��ebr����N�@į��ڇ��'j�>_˼Jx�A��L����;p��\������t@�$���(���1��[n�gw�@Ό�#Fא�s*G\{g��N�r��� ��_E��Ô�a�m���8^��C(�ΞY��ml��P�rOp����Oս[���DiwU�Pu��/��,G4S���t,��5���&�L��U�����wSߺ®�l��jߘ�c�#}��ɕ�7	��˝�da�*:��*�,��0P:��Ճy�u��#V��c`Um��Whˡ�^z�_�z�1��PlRj9$E�@&E.�K�M��[�lx�M�.�:�t�2�����/����#P�� @����|o3�y�6�E�כ���Q}�M�<�n�=𺑇��GfH��q����^�/D9m38Xǫ�a��Nk�.����`3����#���r4#E���z��!�5s�v�3��w�(��xV�4K��\2��[��kB�@�0@�5]����/��*[�^�|}ShB[�C�"��K���:|:;,1�1Ch�� �Ed��"[�,=�BF�?F_��f��Y�5�8��n�6�����a
|$�wk�mG[�'�ݑmN&@�ao,�?yFS}�s����(8�m��PU���Of��e��b2��}�n�U�S/�heYPLJ����ó�F?##�"5��[�h�@�<�-�þ�����~M���:N��P�,�s�<#�l/� 73��f�c蚹���O��7�S^����گ���IU��=�e��+4b��Em�C�<��8G(��M�+�� =³z�~'It>��wL���_Z� b2H��"��x]��g���}0�;#���٤pm�Y)�^Y	����!�J��������Y��
Z����^�=�r���X�p5f���� ���X�I[:h3y�>g�Z�����so�n��68"��J\M���Z���v�����(I��ڀ����o9�H�*�j�2�(t\x�U�Q��VI<�fʅ�>�5�4;��ځ~6r6P\�5�إƖD���&D����t�հ쑔X��ƃ+7k:���<zw�D%	��~�B2Wf�J�=~_.=�~XN�����	IO����3sT,��X�RJ(DOR�Α�QS�Y�0N<��A٘�wﶶ�id�~ǒL#�*���%�G��{�rҶ������j��/9~]���M���"9�q@t��D1-0u�8$�nyץ��W�e��|�Z��V	.H3Sc�V��s����cd~6]K �b �nE�X�]Ȍz/s�϶5��s:��^��% ���E��*8��t����R���d��1`qH8��K�M~|�i�����Q�&e��T���
���g��#,CS����MeI�H"��U�m��c{�W%���g�Eb�P��ՠL� ����Ai!Sa1'��hB�{�#ؠ �2�m)R��j���h�ݜ�iG#�f}]ώ���Gv�.�/ќUqv �{H�x]0��R2�8�����N�V�C�n�@»b�t�R��j^���T��
3�#�i@�`y&7G���$��&kѲP@��4����z�C��e�Փ����.�ɚ�p����z�
*k�%�R�)ꖔR,�E�[�͆l�%F㩯�_�� �"�&��DJ�q���34���B���� �"){M�(h2c�[㜇�m*���phſD$_f�����g��-��6�G��s҅�	��=�y��zk�*Ex�-�Y!cdt|i�0q)KBU��t�QP��W��6ۧJ [���eИ9�?-�?�B�8�(�cB�����GV�ʩ��d����0"�+�����hO:��>$�%`�M?&݅�4Tb	m{���˪,�h|�׍��:9wo4k��y�j�Z��%àCsR17N�W@f3��(�	@�4=1'v˻�x]is4�2:�-1ä�>���RA`$����p�Р~�'E�g�qb��P�]1�;�� �V�UUz�E�W��׽��SL���o��.Dq5����"�������;/��*b���������"4v�5ޞ��c��H~7�&��gnJ"�k����B�� _į�\�̏���9殔���"��pԢ��娊ލ�V�;���7�<A�׀����p��<Ԧ[��Ͼ�3�ͩz  _Q��%��a���"��*�ie��\�3.� ,����(-���-ͫ�p�B�u���2������1B�nl?� ·�"��We�rQ�MO���[�
�������\,��ύ����iK����Bp�fڠ�x�Va?���fu(y�݌�����6}T�9���t:��h����hkr6ޥ`y���rU����'?$�����-ר���Z���)��n�b�z�`�0e�)MCj�LA�[�BY{��;�\J����#� FE�=���4gK�@
����Ep�r
���Zo]�	 �\�$%D:��j6	IO�>�������@g�n���P �����K�N�G���z�O��"��7�S�Co�৛��k��3p�����|���M��D�WN��st��"Hvm�	�AN~[����I�@�Vg����&��%�D�gX������3���'����u�N��S�:=;T�C���[�{x3�����]�{��<C|���M���Z\�ڵ9\HCU�Rp�V�H��`�3h��qb�:���r���"�n�T�������i꒰��� �d�9��m��l~�����c]����m{mb�)p��C;��8�C�KYY悓����놗B�%Z�x�0��t���:\k'��d�]�92��ä-~Z�a�o�"s�p�Z�H�O�)�"��Q7�#��I�ۉXv� ��Cz�P��zVK^�_fH��M�26y���J�
��]�
�٤��J�4�Ӊ��5��
�x��?������a-a�`zV_��p�~$_e�t$VXSlɳTɋ���b��}�nDس������)�P��҆��+R�X�i:8ᬶ�m���B9wq�7o�P�2��#�����_@D܇�T��fێ>�u�s��`��n�gh<�W���󊠸��D��pg�'IH�CѬd�^H*��,��nq݁i?o��J�j�=>BF䮪�ɾY�0�ޒ��d�2T��4ƗD�C��VA�N
(˨4�UBA��^[`��Ņ��;qb���~]=7(���p�=�m�3�VZ��W�g�V�� �D�����VˆԂ0�ىS�Y�	�d-u$�K��9����[] �桋��9q؀�f�Q3N9����H��l��<3�]�%@��A��ij��Xtk0�2RI��Tl�i���u��^5:����,wm�n�n�p�I<^�#%�|���?�ˋ�pofd���� �����>�.���2���L������G���L=dV��cp^�Ӵ-�9&uEη\vl`ƹf�{��RA�|Ioh�',�Y�(�M0\-�*/�s���3z���q��'z��eˇ�gA/	�QGS���]���k��w���8�������y�+�M�c(t
0m��~�c��ϔ+��%��rk�PW�m�/����?!L��,��"18i��Y++��Q�	S>F�mHw(��8��h���(��q��c�������	�j�6泊�z����`�̯�P�0��>+�dAAsi���9E�[u�y8���fQF�>DJ;�߷GC�jj��Hp�����"�Ah�d\m�C�0�㿥ˢu�3�O�R�����K��%M���I�b������`���g"�Y|Xł��U-��!�EM ����O��"���ar�&�)$Ӑ�V>02�h���io��"|���Ё�����M��Fq�)�������\����*U�1	D��?~�TV����p��d�ͬ��
5��_�\�ʜr� ��iXs�����$D�yM�dL?�ZMQ�}TY�yO0���y��|i
3u���!ˇ��,V�/��\X\��N�Fdr�2=yW3����Y���7y�dF�rQnw1�I��O��k��/�@1�V�G�械��Ƃ��&�~W�==a,!sL�O�L��s��w]����m蒕#�5����8����V!:��B3dgZIL�5~(0��Ĺt�������x��./C`'���V���
������ؙ���3�[E�Q�k�yad��1�C����l��]�.fx/��n�lX�5.Ԭ����#{�"b�b_؄�����G��ڈ8�.B���� `�G8�Nn_^�n�ùp�ō��S&���`7�dW��u$r��ކ�����@��	9:;6��㆛�g��y����@[Y#nӦu,���]ҷ���(�ZBS:�����o6<���=pH�E��|9��%!g�+)����ʦ������@C�'|���L�12뤣EHk��z�'��ߍ`�N�1�V1�|6fJ��tT����'s���O���@�ɉ��l���Q�&�>=H�ً�s�k�aL��*��܀��5.t� �������O��> � �);\��N!��@4��+�L�qr�M������o+ %�H�|�P�{uq-U ft�"NI��e�"I��n�9 xl0�,\��S�J�E�(7�i�t�Z ����Y�ӷ��昋�#�?��%d�����C[WyA��"���)6k�8ؖ0�#��O�iSjb�Ѻ��ELs��Ѡ��?���,��9T��MǨ�cѤ� �����ɣ@�������(��|�J��Jiz>�o-�ü�� KI���kt�t"��	��M!���x�w.B)T����g�.p_Cb5��6.QBQv{��rH!"tr`���$��k�S܌K����5w��S�0Um����|��r>_/�z��qz�S���{E�G��J�4���&#�v�x1��-*l]���W�X���1��>-�3�V�!/��C�sTKh�w�V��#��S��0�H|�:�QP=�S��Ae`7������!�d�Do]ϖ��%��<�>4_6�t�^���;�o��+փv�2�*��A@e��9���3�O׾b� �ә>����m�*��;A�wy�� &"���IT�r�|I���Y3!U}1��� ���^Cw��i�(�!^%�c��8,+A��*��	�a|T���|��S�g�eJw��2
�pXk��a �ҐӺx1?�L�@B~�g),��;�G�\�W+v
y��c>+v,$�E�w	!�o�.��0��X#�X�|b/��
����6
���aw�`��j?�9���b4#��2-���J�y��]�G��bp��]�E����'8���*9����Yx�(�W�Kc>��$;k�n"�Q\���~�
�~)_�W|O�L��q�-Y{�X��X� ��Q��h"��M���=t>�*����p03[Iq����n�bpU�[t]l|�VN<����|���q{3v�۸���c�&p�c9������@^�K��ut>Ѵ���aZ��;�b�Z�i
���/�0���P�f�~�j|�*�Z��Àe �(��_�o���PS���q�@�;Ҥ����>ǳ�a&%�w�=��+�."S��q��g�ZQ���x�U��6K�M@%��N`�e�x���A�Mk�2~!������Pos��U����ۙ�3��	���=� y�T�Y=�^��=&"3����d@[��� �rIv�mHէ�U�u\Z�%��s�M�%��ln--<�kd�l�$�����Dw������}_�I�(w���o�6vP����A��If���mw=��.:�5-`f���Vm�()�I6�՛��瞶�^�A�۲��ҕ�4I��M�)C�^��K���c >cdk3�	^�*&�y`����ҙ����� ��.���dJ+�A���Q�ܜ��b� ����0�>S�4G��
��w���fZ��q��1	�돆��u�{�w��R�
n�O�r��s�y�A����> ���.�0�J�F�N�	W*3�2�(682(���yV��<_jo�K(������0J�\`�A��7��֠��i݆%] 8���"�Y)5�3�fl�>j�Z.puug���zE��99�H[I+� �;	d�U�*�3��Aj՞���+q�R�&%<�����j�	��W߀v���_�Rt�fB�;"���'�yb5�.Յ(y��F�Qv���y��˂Ey��\�,�l��8�`-�(�W �9La٠�)���/liAe�w�k;�� �Z��"���Uzy&�r&�����qs�P��������y���s �ty	�ӈ1is]s��d�d���O�;�ͩL{�X�ɝ����@7dGz{M���wMC�Λ2G�\�H�"��g���s#kܪq�I��$,ق��2���Mr�M�N���bM0�� �/}�Z,�f�F_ٿ��Fo�k��5�cJ�r3�6/(@#P���Uk�GLv]�%R�Ҋw��M�~9E[�s�b��z3N!�g7����ܷE�4`�MM��盹�,�	�d���n�Zc����z0��j+nQ�^���/�`�J�N�>�I"]���0څQ���>��A��P?�I;���r� NX�p륌k����X��`�-��i��;)R+�ĥ�.,� �gSkW�f��ɕ��\|?�cv`*�#ˈ3Jh=u�x�=u4	�!c�/�c���,H��
|��`�1P��2q��U3��z>��3:���(S�c���f�����܀�[�����9�r�`��+�&����XI ��e8��y�0�>l���V��	�l���#�x~/(R}��÷��p��a����y���S���ʧY�wT$���00��X��ب��%d<N%�[�����M��^��A��檰F �NP�\�S,0�� Ԋ��I�ݒ<��>����]��#]� �~(�Y�9����U�U��<��%C
t�%й��J�3�t3��׆yU���ȿ����a�&һO�ax8��