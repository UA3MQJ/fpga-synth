��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�
���B�+�3�I���?��n{�w���Y�2�XaUX�f�>��X���tx:cJĪ��\�ɿ*��4�����I,JA�S��U���~o��(<�
���O�"h�f��EI����.��u�e"�����y�~N�Zl���wq�4��q����G��;�X'_`�_�
�)�?L�����
��yN*���e�k.Z���s��
do���+�Ct��׺@��wۼ��c%6&U�n�j�l�q���2�6�y�;w����,��Z0[�k&ސzz��*T�2�-�ѹktuCQGl���egQ��`�gex������bc$1q��_�
{���v�T9P���'�1����'�O��<��t��Aɳ"�b����^?���!�Ij�W-Q"W�OA��3�G
�P�t,��l ��Jʿ���9� )7�'Y��;U3=�j.Hdo�.�F�z�E��k��l�QlN��������ؑ���0cUE�����p��st�|�������?e�ϋ��O�y|��A��d�r��9�Kh�C�	.p\�
�å�.���aԧ����7��@���>���>9Q�b�DX�W��䏯��C���ځ��R��V��7
&C���:q��1S��݊��#,b�*�2g��̒��a0wSD0,�uE�C�`��j��H��@��Ϥ�}�.�%a&����w ��� #�j��ҳux��������n�����3���t��m|�r��9C�J����
i��ֶ0krt��� Y~��~X�a���0M�v<�9���r�V����rl��c�BU����������%R�
[Ђ����X
�Bsf�z�a�|gM�uC�c�� ��hc�]�#���d��Uwa��΀\�� Lx���j�k1
����ۿ(v��	S�	bp�$���"��a>$����В�K������V9�^�6�:�PA�����^�S0448��;�w���#	���|����Ƕ�л�&��S!u���D�1D��ث�};>��^vk���ג/r����L�#�j��p���� 8���\��V��d�����Ƹ���
b>b�6���H�H�"�lS!9��y�X��a���;[~xi�s5���	����{\�L�z4�jXC�#����@^(̭��9s�{��{̚����b�.����GYL_g�2Ӏ8�qf�0���益Ex�b�yث~�$�q�h9	�$^����T5�v?V4#�x�yf
����E���DXNN3*q�gbˣ��<)-#c��Ͻ��d�ߌc����#`��QT\}��EJ�a��TKU+j���U���r��z۳�)E�t<%#u�
$D����YJMa��V�Ҍ�v�v��������fD�{6�[�� pn��.&̚Uۉ:�2��Ǽ
"�2Y���B�Q\m�`,餌�e�Rw��D�z@�DXe�Y��qʺ�������;���qhDo��;	�o�{���f���Q��$����C�w��T�8��Η��}���v,�%�-T�P��
=C�[�'\=z�BeQ;����Z�'�����A���p�w0���1��q�b��<�fi�y��y��N.�@&v~�<u�f���ϊLjBj}>�{s��0o�JK<$
M&�)w�=K�2�8Y�lo�OG^EZ��6���~i��DHY���^z	Ә�����B�א�?�ԕF�ݿv�sz��.Sۀވ�Ҩ�����H ��|�E�Y;�{4�xu��2�Y�
֫�Cܳ���tPP�~*+JN9:�W%o.�C� ���T�e7�LXr�OS�*���%Y��s�����k��^��I�	�����PFz�gr���թ@&H�\�Waȹ���@��ό~�3C��]kb��\#K�ވ�DS"�ak�7���@V���ޔ1�@�A���\�B ��d���9���֠D���}Q�뿐WC�8��
������64a��G.�h�P�b,�F�jR�b&"��_1�d��Z���(�nA!�&��4ҏ�k8�O�A3�T�u�A�B-.o3氃�(��?�{�	�e#j ��g�B���G_�]FG0�S�Ȁ.�7F�9i����7$'}��_NTlH�!*��Y\(���]N��#�u-x"��ۅ��Vu�6���Jz���h�`�UK��w�!+�~Ki9i%���N���"�+��
)��6��͏�aT! �!�S�Li��Շ��H��R0�k�[OK���9��`A���q���;,�((��O����@�"����<P����A�MRx8��w����ӂ��̭�O�Q��M
�Y�R;�Tx��G"�����4�, ��1���@ �m@m�(d�q 
_�i�9��T�3���ڦ��t�+�����+9��|�`�Z`}K�{�UI){���Wg�(��+�:��)� ��h�nu���I�J�L�
�ⵛg�h#H�T��tn��\i���|"��m�6aNfyY��M����DB
:�n�cpӬ�h�4L��D�Nd�(�y<Q>�FAI�4@�[��4�:�~�A6����9�hᝠuKB��h1�W3��<siƭ�-��^�8yb�,���4g2�������T*.ж��5=�	V��l�/��8>���}���'MDf�\� �wr���KMt�JH�&�t~�aO��4y����l��MKe����N�S:G*��Έ�Z��e^4��^p���c���3�1:�Ւo� s=�y�l���a>Bi������.g"��d�i�[*�$<�6�����Z꬐��w����%ő�/�SƂa�¯G��!�(���B�0qw��u|Jp7h�Ȩ���F-���9�f�k�]��)��M?�f��:
Z���c��@����D�&Ѭ��L�goj��:�]�5/x
���w��g^S�����٤D|�A�i�rK��XM�)Ǒ>��'p�v�����73�{�F򩛯�v�S ��ty�Q���_�3�����a<Q�����Ԭ=����78��N�����	�`�C;�����=�z-����v��̃4����DժW��ܺN�8�p� 5+��'�*7����_4�{��q/�R�=U[��L}}����yi^�j�SS��*q!�܏�]�n�`	�o��q�B�6�`�e5}w�J4y�)$�1k�w%ot7b���yP��{��� y��V��(�nnPl�j����{����4�6\E�0|:	�j�!��)���Un�+�y`����궵CA{fLP�i��Ӝ�ZL�wy{����'1�R��0�k��-l�c�>�S] ����@N�6�2g7q�Ih�N��"�Y��kS��� b43��:q���Ԝ�<�ͥ��~����x���QS
}��!�tx���qǘ;Q�{{������%y�}���i�
�����Ï ��	���&;�6�Zh'DUF���t���h�~Ǵ[HV �,���]�ui×i�3�ſ���8x��nqg9��ldݗ���@�v���%����������k��Fl�[�qIez	B� �V?B �4�k]����:�C`\V�Z,��E�u�R��2�y�������إ�h9�a#˗Z>s���K�ز�Z�� �H������9.M��&��9�(��\s�=+m�4�;oOR�R�AF�;�s����[+k�a�0�]׾��h���j����|�Q�U�DV����o8B�u$�أ��-��]����c�2��=&��y&7(��>�^t������qސ���q����|�T��� j8�.f8�{�
-d�m��
�|�H�
�(ׇc0���al��:�F3&��#~o�'V��Z����{����:���,��PF�I�X��B�!-�b�l�
B�Y�ۣ٢vN��D�V����L4�R�� ��"�ȿ�l�J}m>LGW6�%�H23�j�
�K��a͹����"&�o-2_ڬ��̇��z�iu9�]au#�JY�+nZ��Ғ�հH�(=C(
b�R�h:qm�A�]&�$I	 *�������l��>�]�����i�}�7=�	f!g��JO��=��U��	Wp*ǚd)a�QǛ#-xt��o/*�1�J뷹�ԫ��i�/���dk՘�����e�|����>x��F/�z�ч��@"�2R�H�����~��m���@+eԈJ��of��o:�Sr8���rz�W:�겸%8���Qp����f��%��-�݌TX{Hm��L�S�(�7������v��;D��=&��T�o!�5];k�~ש����d���t,�Ȋ7wd����،���/Y���ܚuNF�s�b^K�$������t˧��w/�!�嬝W�&�R8Ƶ��-�K52x�>	X�0�|vv���E��g����I�B뗵wT谢�Q)�B]����b2Y�l�#2Ѥ���Ժ�AWD��\Y�
V3B��32��]��������%�yy 3��~jZ��#t�f�9{x͒�f�D�����j�3��y����˒Ct}B����A��jp{nW��QPѩ��0�_�6Nm4;"XWk�Э٨9���՞�#wo��G ?��Fj�+��%#�`��;;Plѳ�Kw���0�y�;�f�Oe\Z�Y%O�<��	b���F����3�ڷ2���/�5�&7_�h��0fg����s ��d.��ٸ��8��t)���3������;��z{��ω�C�ŰV�����L ���|��(���v�.d�X~�k-��z��:��<�{Rː<ezc��L䠥8��9�����V�r�hm���;�@��S�K����h�מ���{�[����m��c�iT���`�Rzo,QB�hn��ڵ�[wt�X��|����y�K�7��A?]M9�Vgq��hg�
3����]��:�DNZ���2e:f'D��R�6FY0iv����~H_����G<�l�c�V�x�)���~2�K�dKA�
�<�}�AB������C魽�>��=�0�:��d"��"�),�Y� ��o�B�
1G@��U�?b;;�$��U�n8� �f<y8�5L吗;	�_{��xh���l�����k�ڿNfS�a'U＃�XL��mtQ���5���5'�F4�.jk���h8�|K�M���Ml�E�mW ��Q�w�\�d�Ԗ�]S�;�l��\I�g��;�v��F��eh�����$�I��)�g;�`?��'׏'���%��שr��t�z�;��ZW���+w� .e�'�l�,V9�%*����9�^3%�Q;�쟠u���;_�v��?)?�jY�`�	�_"�
�]��L��z~��G5�x���``J�J@2�|��R��cy3DC:\�K#�13'�Y�B��2�����&z�(�N �+Y���I`f��6�n�� I�֥qF��u��K�n)
�}� I`�Ѫ�SP�f��q|â�Z�>V��tȠ�A� �Y���D��֩ �Ci8����Pv�kQy^�3����C���꛿�MY��@�8� �f�L��FY�`�&�������{?A��*@�^����[���2���c|�P�]�#'XL�.Cq�߾_�zį�Ѓ�p���丬�1�gO�=z­g��ʆg��ߖ�t%����
�n��aH����p�c8����8����d0�A�Ǝ(�?E�c�U�*q���l4�P�O�@[!N�ȡJq>�C��"�7\�SnK��q��F��NT���kjn�`o��Ԅ-�M]���K+<�Y��R�����RR�N�q�61�9ט �Þܪ
��8�����NoWI�$�����G	��^����+�Z5
V�d��=˕��Rd�B�K��59ͭ��0�)�����������W ��T(?��T�!�)�n�:墷�ƼiQo���l��i���4�m/Fю�1� h^�)��W`���ZNiC9��"�ڃռ���Lr�?�+	\32|�v����r9Ȋz}S���o�����h8TB��ҹ�s[�U�_�a�� ��\�X�Ŕ�n'�%�d*J5YU] �k�*��՗kD"ςbi�6���K��$�y|)�7�om��<�0u�|kQ���̝�h��!R�@sZ��6:�������n���� �ǒ�7�`����a�TTLRRqr�b ��V�*n�m<�I]vY�=l��OY���@��m��Nu���'d��O(]g��ݗ�r.�j�:���+ap�YޥB�RH�� �N��^X�l�w@��W�������eq+�^C�?ȩ�:ߢy^�Φe�T_����DK�N+^��ec�� �s������"����.��a��>�T`��H�����Dl26����к�/P�m���P�@x;	�# #�]���P�P�gd��r��q��ː��L����)?�cM�M�(wV��a���Bd�.3jo�t4&�d��[j0K��~�*ˈ�'�@��}�Y2i|"f��aփZS��a�;��{�BIY��4��يVf~��?�9�j�h��%�k	�h�
3�}밭i���c��������o����;v�_gZ��l���U�b.��--�W� �ށ���l�I�ڹ4.�y�W�m
�2�\��r]�[��x�S"��+�Dv�������~�Y��O�n��BLs
�����=���p>�RHO3,�����J�Ưp���ZT����;��7.M��Q���3��W��*��i�����T����Q[�[\wOp�z��&,������k;��+[�s��`krR����%��^ʬ�@|�Q҂�R���^�C�~%/�c�l��$�U(|��u(��X��-5�����?��&hB��y�9�5��QQu�L*��7��l��n���b�Z�TJ���
	�R� �m	%p}���B$��\�*)�#��(��"��Y�P��x��6��KA8 	K�m���ů�� )	�'��Z^ɫ]��s+;�*%*���"))�?�#�#ϱ�ݫ\��6C�C��t(+�6�y��v���J�5y�5�ٽ9L�ZB��*�O"*�)ֆk�ةq�?�g5eܝ��p�3�ӭ,&z�q ��ȸ�e��IB{�gRVzd���01}�i���@�@�%��pPu�d�2ix��c쯭�⇗z?S�p�r-�u�Nj�E�"��(�r�io�B�:���O�wG�
�eO�6YL���#W��ʯO:d����'1A$�f�;<�� �����fE����71e�C�>����('v2.!N��^%�\��zyL�h��j�Rܼ$��;�k�o�Gaq���e�|S���6mٿ�%�)�&�"�u�u�<-J*�P#�Y-�t:Ƃ�}8Ki��VǮ�#��Z�5ai��Yx0�^�5TA��������~}L:
�a5 �j�O���ٜ�z�-L/�nӁf����B�d��:� �����v{y.�����{���6��ڛ��#�)�U����#�0�OҎJ�]�]�ߔk�8��`	�2�ELkE���:apw�I[����C����Pr)�����Zuv��
*�]8]K�h�x��
<�p�?]��B��������l%z�GCB�G u�-ȍ�DX���h�)���Ǯf�:��P�����k��/��pF>�[�c>ϣ�^�2��.�p�g�A��*p}�/�R��70���\;9p�=�8�%(����cV�m�r�2��#!<��T����^Q���;z�%$��L�2� �M	��gafqmds��6X8P$�p�gX���dś=:Ɨ5JH�<Mt�]�TxA3�(�cP U�pQ���� ���W��Mr�0��Bc� K�i�xQ�����'�b�|B�{]�
�&�mޢ5�ݙ/�T�V�H�B<=9���(��z��{�$!$rg��Z��+�8޾,�^zKe��~M�	c��մb����1�k�h=�k�}O�g�<�������yIi?�b��d��T�ɕJeu3��F�֌�����[�4+R��e&v7Ŏ�E�P;�H��Õ
�<���U�
�[׌c�աݴ.v	
�^����4<� �M�Ek�A���7�B���˓'d�]۷�I�9c�S�k�����퉿4��9�Sl5v�|ו�o`�#/K�Z��� TA�5�V���/)[��E��C�lK��)�E_	�׏���s�P��������9X%gY��,h�"�]��Bi��{��w�Z[F���l.Ff�fD�N��qo¾Z�9@%L�ln��a���P������T������ 9�68J�F
j�o��/�\ʡ��K!&ފ�ޥ������PiX�Q��F����Ÿ�Δ�w��M8	� �NT�4�����N�#o�IH�t���^j��r9��T��*�Fxe���ٝ���h�vFǎ���V�:`+���<[�=)Pӈм�T���pؿ�,�O�9%$u7�ʄ?��1�0�t���B%r�N�^6L��M���Ke����6����1^�6$)�p
/�L��^����T��}_��?��P���5a���+9�5DNiJ�g�q�gE�=0U��C�s���37�
�
u��h�H�=������H�����D��.	K�`��߱� �S<f¨(9��ժd�{���KW���V��m��F����.��s;���@+;L_�ʽ,�F��C��~R��4���8S?�!���']H�$P�2��q Ec�'��18���rY�O9po�9	��y+L�������S�L)�K�\u��P��l=��M���0�5O�ު��i��RK�"ߺ�������)+����XB�^��`�#�d�+���s���:ҥ��E�_����~_������P믂VT��3�������k�P�߷��Ďߐ�i��/�^�Y�"�sG9\.��%L�#{���Y�n���8o���`�o�ǭ��!�E\���9ѵǲ����Nkd��z��c-ni�C�I�a�(��w�A�r{lls
� ŝ��w%�Q�p��}�ϕ��d[��v��@�/d$ �J�BMXr���E��]���LF�sgx�0������o�A�ԝM-F�l��;���s"��{�o�`.����ܰ�X�oC������9 ���8�I��[vi�g�T�-�E������|��B���nW޻�����V~%�?��%13Q��ͣE��H�T�+��"��T�o*Ǣ�7 b(�M�:r3jj����B^�X;ݍͰr��1��N�� ��T��o �����	�ā
�P�k�99*����G4�i��9U�	��c:Z�;��D����������з}��EU����׈�oMQ�~���UT������~��y.�#����k� ��H���K<E�sf׊' �M�:�N�P�A��Կ?0����z��N������wJ �,�J*���᱿���,0�*��0�Dd�D�19�OY<t%��	u���?6�b'���\i�T�,��f펝�E��Y��� N�����@��x�{s����$c��9^Y�6�p�u|�^c�MV7��1.��X<�k,������4�����p8х���@483��Ĺ$e`����%-DZ]��O��Y��CŽX ��ğ�ޮ\�3�
�ى���.��6O�E!9�sDi�e#b�0í3�r�W:�E��"�&���CA�6�|��*�90����Mr��M���8o�2�kq\�_v�ڐ���¾�"���yeU`��)*��.����B\�w�ﱔ�4�:éQ�B"�}�T��XT�ß���64zټ��?��s��J�}�k`�,���f߰��(�^s׿����B�J���"X�>:����E��Gs���}y��8}ˮlfe�o�h@����U�Ù�%�=A`�m+�2=e��@ p���?�=��P�]��_S3쒘#��T媊�<��jD�R��!���]�����I=n!ߓ��v��$yNϐ�d�3 A�:R�N��t%��{�P,!m��ľ�ޒ���-n���y"��s}�C����ZI����!�U�/e�Gz��L{nvZ��v_MH8�ތ`:z��%��f���,�f���y���$� ����ǔk~U�1W�PELU�"���ĵ����E�ح�.�~zq�8j{��l�Tx�Kq�]��&�_�6"����8gx����(��<.u����������߮��3h�h�qWo��% t�R	9s��쭛���1B]1��RFuJ�0@��y����f�IZ�A�h��.&Tn��7)�:���%�!o��� �B�����5�Ő��'ٰO����_+h@����H��{2S���p;���dz���f�#�6���;��,�ð��½�jo��S��n��X������Su�G�&M�U!a��M�?���,�H_��D�Xۛa�����f��Heij����RL*�P 	p!�,O,��df�@##CN����3�2:<<[�O���&���j�]�~4���[�R�ø>�A�����d0�B^py�@ߘL=��N)M6T�����TI�{�=J��ɞ�rV��x��T���K2��	����-�2�,S1��@���s�9Z��b�*:��o�bJ�x��Ée�I��􆁚NO'U<Lo�`�]�o$�i
TlK������519x{R���ib|�~I����2%oᯐ�䠙�Bv�x��#�ׂ�����k<���ɜ�'�{�l�abJ�u�ݟ�yh;	��ر�V���N�p�ɠ��;��.�	�T翀�� �
.yO���E�!ɚ���_��!f�����(]�A���Xr�&��2��w6,M𿷐�s���RY�~���L�� jj���=t�V)LW��5��F{a�1=���6jB��+��-�q*�7IC�<���E�Icȿ���y�f�}:2��{A=p�K���Lc�݌�X����F�F��s;������VL��v�G��\�1	!�lO	7M�Ⱥ,��w�����ʏ͙L�\�	 N��;���:�J�s����T�Z��rj��5 ��(�U�
��Fd�s��ϰd� !B�h��-�wʳ�0�Jc��=&�gB�h�M���9�� �9�c���c	���#��9�1%��̲������ a<1Tue���'�t�ȖA]?#*E,2��tH�B�;mᯃ.����ڭC�x4��U����^��$`mS�kG�y�F���w�B��h`���H��UW#0�N�Qk���ra���n"�:�jc���<�?E��H��]���0~�5�=_�}i8OE}/����.M_��_6< �S��Z�1`�P �i�*�̕���c/ �r$��s�$�jխ��M�QƖ��-�arKRM���P�AX��d���.�N��X4��������m|��c�:���J�ɏ��XM���}�4tG���'�&X���4�ּb�dj���q~��w��mƕ�8����[;#��V���ʬ�.��3���#�?�<�b����՚rP�r~v`X��0�j�I0����Qc�����NzO�Gm� L-*����|}⫲�c[_�l�11jG�&�Ǖ)J7R��?k��Mͪ6qWv�E��� I��h�L���L�t����À���������j�c8JA[+W�b<��p9o��Ԕ�qyT�Y�ktx���@�(%A��N;u%�� ���8�zM}.8q�q�(�w�'JW�q��Z�Zg!m��3��O7��f�X߶.�)� CԤhdʨO�]�F��B���
�N' �"�_�F��a@���*h�S�<-��_��CU��m��V���P�*Y�z�P���T0�*W��b����[�җ­�~U&LgfSC��%���'w�I�䶑�g���S�$�1���?̋��٥�ɑ脆�D(��xkٱJ0���s���$�s�	��Â�0�ҏ�����:.���aj�H��&K�&d��/m�9P�(A���[�FK���á���n1Ϣ�(5���TyBm�շ��sb�sb5T�T@�{�d��?�ք���H�=�ّ�8,���ϭ�kV��k!#p��3P}S��/_��L<q'�,�3�dt�VP3���	��E�ܻ�b��4��w,+�6���$A�Ch��_lh�ʕ��a�#yV��z-gޯea
��*"�w+����Q/��G9?�};5����n�|�<!G�"Ih���/��aU/a�e��x�,{P7p���9�i��8f*IJO��D��g�{p�ɭc����5t� #Ԇ�ػgm���%������W۰|����ٔM�.��>�0	?a|�(��$ȥ�Lk����L���}���� H�uD���>�X��*F�-�x�/)OXYt����WN΁�QNâxu:�vْ���g3ob?>I7%X��.���wjx*��B�*�ф�� ��
������g��	<���X��;c]*� k�9�Bt�&�r�XRG�$���c*	�.vs�4�l��z�����hm ��x��ލ�*m���-���ˏV�u7�M�C���QbaaA)�6�:?�M�ce֤����-v��}t�,P�ac53�c'����D�o�Qÿ���nW��Tjd
FF���	y^b('�`2�~-?m��x�<�!i�]DO�dc�L��G�g��U��K��L^����:{��b�W���2&(pսTH����<5�x���}�슺�x�7��س�g�Tm�S����Q�<w��9�:�ضM�{r-F��Qbh6�͟��Xm`�^��j�!_SA�$ظy�4�� x������Q.����QS�u��c��,�|���R�	(^+I���|go�QTDo[�b4��kʴ�- _D�Wb���'"�G�Z���'}9~	v	BQ]6���@��^���ŝ	�BbقP���-6�r;�M7G0%k��`���3�!�X�i��]���4�K�4�^���|�����tr��%)y�p|��y�Ũ�G~�H�Ą¶�,K`$?W �vvDM}���*���4x��,`�Q�L��W)'����\��JO/blB3�[�}��t��۠Fi�hi7?]��Og�%K�~n������'a��th��2fZ�w��[Rr(����;p��{��fZ�߽��a���j(a'&���*�se{"4Ӻmsר͇����S�i׻�fL{$ЬҐ������`74�e�!��zb�����ʣl*��d�6�a^�%W�V�4���k*Y�X'��;=�^8�;�^�r��F����r�ʄ$�b�KBx!.��Pi5���X�����7�{�g�{������~qə�Px[��׭mF��3:H{�"/x���@E-�m�a�9;�al�<�/���h�x|�WE�_h��ѕ�W������,5�C��!��Ӓ˧Ƹ�,��ċf�[e��&���?ي�B)�������BWX+�CU�ƪ�ķE4g�:7��L>�	\aF��ǝ��Z��@Y�;��ʵ��g�[@��p�}`ޮ�e9sF��P��JY�
�n�C��7�$�S��2ep��ȅ�������6�
i�.͕@�� ��=�l�"﷬���<G�}q$�K��{�H��Zf�(i����E=���|�J=+��Ť2Gb��1$hS���g^F�eV1��L����}�)`�b͢_���G=���Hx,(��FFۤ5�w�8�1vP�����@СT���Q��ī@@�>�Xp�kխ�\��9э��+V�af���=?�WI�A&#�.ƕ�9�w5��ZE����m8�̄�⟔3q*���OIc_�OAϪ�&j#^uR�DYLj�%XK�O�5](�S!5̅���,��g,��]�*��pYZ�G����"�{ſ��cy��cs���%�VJ%�r������*��U_�.ղ*Z�im����Ԏ�E�'���4�G@r����(4��E�(�a�ݎ��z?��@3.�����q���5t�B�,Z��P���e]/�j��%w @f��p��K�,NS�߼���� h�k��O�<<�`��tp�<�8���2����O��Σ%P������IX���[ӟ�EJO�ok��K�"BV�����O�!�*�4�k�_�[���`<c77;�������م���DQ�re������E{m�ϣ];X��38��7:E�bO�Cvk��9��n��o�wgwo,ra����iU����ە��n�D��?f*�u$ܞp��Dӕ��(%��Y����C[��	�!3W)H%��c_��ǯ�5I������L���HtEߗԞA����B�����M��>QKW��W�ŪH�ү'S��|\�e��T�lD�f���e%{	3bN�� v2�y���?�N�8�C�#��+���}���V�hav3Z�u��Q7�:P�ub7OJ��Rzs��^x1�!c{@6O"�u����S�2� )6\m4{_�	�Ş���G�u[�f��x�t؈��#	x��y��)LZR��Cp�7t�Y��QK���� ����?�2����u�l�X���<"�}Xx��蠉�wX����hz�:�M�-L��mUSŻ��tV�&�sw�d�r���9��|7��!���wM q��=V��DgRG]ػ�@[{l<�}���N��l�e!|��]a5�����"����N�z�&`-�'Wa���	5ɪ��p���h���zw��Tz12��m�S�%�
���.�yeЁ�{[L�r����ؘJ�Ԫ��x3��*�f�U�f�E��4RO`2FD�$�Y��˼�rT��0f�s���}�	������N20���Sjr��� �8̀(/��z�o|�ރy3ǖu�CMn�,5E��\���8�ot�L���e<A�a�k�� :mK&���9k��$_`�P�C�݀�1�-3�Hm��r�M_��s�Q%
�ڠ���ZTrOX�r�VsLއJŅ\t8r���j�'�e|Y�U�Ρt�`k���Z�[V�UY���͸o��Eʴ.a��9����U���9:��T������b�F��t�oWd�ɱx
�|\�IW���S�c���;��v�o������W�^0�0\�٥��,j�B��3�;���U���]�f�$�+V&�Q{�f��܆����:���Q]�N��u�^*Hݻ]���4�Dݐ�J"��I_��2G34ԣJ-�wmw�[�,Zw���8U�w�!1�-BU'��&��4�EBO��M��K^f~���s��A̻d8^��}u�E�dC�����"k��B�	 <�&I�YM�?#�x�^�sޘw���%#1WrYp�H��ɞq�� �2uVt�fovc��V\c	G�L0h�8��hM�,���ă�V1�U��� e���@&�
4[����Q�q�V������l�+�P���֯�a	����H��9"�[��~;������&��h�_`��f��G�rbp�ַ�n�o:��R���ηa��t:�{zV<�P�9�
\���3�%�͌��?��Bq�)X���:�����/b)�ǜ�j��w,���G�%���X�����n��;��^�^�ѿ|�a��O��O��Ǩ�����0�#&?Ј��Iؒ@l4N���j��}���V~���^�beNnF�A1l��C�o��$�;�q�&��?Ѵ���p���T�U,�`��� &pŽ0/<�v��*����Ų�y��M۸�!��W�y,�#	��0XxH�)�X��z-����|>�i���4Ǣ��.U����*H��DF^8ʗμ66B�6��Z㮫uZ��=�� �����&)�R���r�&K_�>S��W��Ezj�d�kKkE�Oe�����vc�`Ct'f�D:p2�V��E`ܘl�=���`Qo~��"l�/_=�REK���q�L��1Cӽ{�Q�:��8 �0B#�bg��uO��G�?���+�x�?�w�]��G���%�S~�tg*�C?H�gz	���ꨡ���(&a�2v�$ �I�qШ��ǭX�0�,A�\��	����׺b�+;?3]Y������y�lUz;��o��� }����a��R�5�9�v:���fk"k��(�o���󇠢-�߫TH����zi�y3� ���K�B8�6n��G&��3 �cfj�<�ko�7�l�P@3ķ{�%yu+_�R���(P�YT����$�-	!�?)�:_��&W�@�͢�����]�7p���]�V�g��o9�I��MM�� 6� �$��{�9<�NoF�B� =h�rc�@����3F�H̶�ك7�w�-�2��ou�7*��Q�^�#�;��х�}&��oߡ,�b��_���`�;��X?-���wObS�'���n���w�E����Ɍ�)���ȟt��n<�[uS�������i_�8y����3�9a��i��<1��``�	B�+R��2
�#��f7\^�S'��\4YLiU܋�\���J#W�m��J�ͫ��
�������1��Qx!����*�đr�H"fc�����ζ+wO佣���.�S��Z�Vpp�'�#�GD�3�V���ܨe~eak�7�/�M~A�
��h87�)9e���S*牔6~iYW44�%��z	d�]�{���������`$"��S"r�����h�e�~��
8�+1u��#H�U�H����HjI��!H����_+�B�-�����b�=L�N=N�E��јbZ��tr�Xk2e�?�!<{��-8z���uO7[�(���'��p~��2�"��^kSG�\��A�M�*�Q�xF'�fdi}X��?��m8n!�ȓ��^Y������k��[�m�ʄ�Ґ��|�L��`4aMY����&�}��˽�)Ve�"��Ǖ@��Ba�㦛 ��k�_pf����7�#�t�����M?�`�YY��`@��xw_<(��%�`_��+��{�0-�7�`q
l�9��I���L����\z��ٟ��3��;�8و=��"����ݿ�S����ܞ��`���������+�P�[��o��qK�ﳪ?�]	�z��­,Փ¤
+��jy���n:�
�6�\ơ8���Q#�Iͥ!������H��ky���+��lЌ���(�+��8�,y)L�N	����{4���h�	�/c��lg��F��ɫ}$!/포7��|�F����]o�j���BלB���m`/�y�E�QV��2/_@X\'_"@�\���$:���ޑ�B��(�]h8����xxJeGm�NX���e�*��~�M����U7V�	* [��j�2g��Y����桪� +sP��9�(i�J�rVV,i�z;�.�`iH���
-%�b���I�#��?����h��r�J{�ǈ9O�T�"�¹_���	[~��2p�:p;D�t���%�؉V]�i"�� �`��q�|�ސ�,b�Gن�����A=v�9VqxY'?l�K��nV�l^ln98��t�08h���X?��hֲ�?�:�<�ݓ�飺��1��i�����Y�ɦ؃���������a,D̴�!	AzH�WB����� 
�1�a
mV^XU�k�|0L)�$�UD�gS��?h<d��I�*5�2�!�V>�)y\;�}��o��s4�`�V%��j,~��oӏi�1z`���M������tA�g��/ʛᠤ�C`fϘ�5m�� �PO]���jܶ����5Ƨ��Ej"��g���g�g2�¡S���Ã�rN�ty��= Ay M�It&���LĐ=F��м��:,K�t��3N�N�3�*3�9����*�HkJ4�VUAͨ��z@i-������s�����7V#��}�ڂfH��Lb��=:[K���8�?aj�Hρ	���?�GB$�����Pjs��u��Z�R�ȏ�3u�;�.�6d�p=ʚ5�/+����i7�h�o�=,}2���8{�K���7O���ebT���j`�N�n����n�z�ȏSߠ�`�w���O�	{lx�����"�����Ye���eY�9�?ִ��gJ�J-�9��~�z��b��[]�ܰ+ϵ���VR�ݡ#ǁ:'�&gh��x���h�#KN��g�~���n��ѳ�Z�x��j5w�HX_Zv��t3՝J���X?��FՉ���<�z5��N/��y���x��-9�	[q#/x>����#��<�&�܇��4PA�7��d��_�o<W=V����Q�2�Ӳ�	fċ��~�	v�Y�����X��'�z�����w/E��"������׻��`�h cN�����^7w�Z�ȣaH9��H#�0ԞT�{�-� �5`Π�Wϟ4��ays7����ZP-;�:����A��	�u&�H�9v�B����gR5��$�~�Oa��4���{����ȏ��?H���Vc�U��kߢvK%%��=S���j�ư��
4g�F�oG�˓@p�����I�~�m�H�P��8�T8��Y���iD3 H��j��Ao+���^6�w�B�od/��I?���O�*J��̚��S�3{�j���J�vF�zE�}���>������b$f�8B��4� ��ܰ+�n�PW�`�l&J�
ԍ�h�|�� `�(���4���X����Ta}��v��R�&�n��8�ESw�7J��H`L
un��h���/9����.��	�A�!5�.�qaGD��F^�`	)�l��VIkU��υE�� 	[��˛�"�%�4H1��1Ϲ"��h_=C;����!|7)t��ް8<��/
���Ҿ�o�M�������.�H}����B��nqvE��P��lIP���\�ʄLr>z/��6v��)�#�-g��V��@60<~[y�7s?�8��f�1���ûZ-�nܿV��n�z�P�!<���t5?�����3Y��2��5 ��ó��V��zx�����:�E_Nx�؛.v���^�=G~%K{�,�I���M�Ԫ�0P������|��17����kT,�Gxc �TO���#XX�&m#��)�����vƂ ���Y��	v0�{L��d��V2�rC��'Ax����;[ۙ�, ��L�]�$��*͛K�TS~��G��R��$���6utB2�C<hroy��up�O��<�ݦ�6
�8�7Œ��`n���i	
2�}>�c��>�9'��s֍�W,6��P��K.�.<y(�Z�P�����ę�'أ��Eӣ��*�P�aH����f��1č�$D�~B�e���&~vR}N�;�]~�J�NH�h�M�&�����|NՏ���d��?���k�FG���Y��Ԑ$'a��5��K��H�ꈂd�6[��� ���sm��_�=E,��Hej�7O��,Ɏ74
6Nmek����5�˺�X�a��w	��؊c����}���h��Ua*}cg�l�=-0�_�4��&�Y��q^su܅�#�RYB
x���(Y�ŝ@���4���o/��8�Z�.$�oa����zs&�&(���$���MP�y�Bf���,PO��>R{��_-y%kv��|h���~ɿ,π��T�^��?���ݲ�W�Qy8��]&�+���~Q������﨧T�U��#@1��'(]��]�jE�Ê�8ݕ rt*4[CU�W&N��T�9��I��:��#��3�'�ے,O�zH�ɚ������Ik����ֶ��d�؞=f����{/`!z�Y��>�.�s�t�+҃�����-A��`β*��p$�z&��yp�MR�=���x����������.G�+M�|�:�OFW�f}@�C���Q?�l�����L��Vg5+�^L����%�.�� f!�<�X�N͒�	�8�E#s��v�G��0k�m'�N4][*�7�S�1�9"R��(�O~,�i�� �}��jp[�]Q��
6M��[
jόl��k������7���_���>��U3��ԺL��jB*]��;-�V�V����38�(�����Pw����ٚ�1�@�`�nj�TOZ�`;�r���4ݓ�!���2Y��@kP̰8wE��hO��_V-���yRj���Q	LiP������B u�'�z\*=x��=5z��'�jQ+���ֶÇ$�)����z�Wm6����B`���p�!����p�ҷ�&�)���8E0�qv \���@�}G�Q�9�G�<e?�C�7����M���!��ϟ��D9�u	��4���P��xp� �#��,}��s!��������UYf'�K	�
�G�vj��8Gfo��]|f{��|�3� b[���x��H8�.��֧�A?��2(Q�=Z��7�- I�\pO�i�zNTa7��\�3%�r����V�Z/B�Ƹe�ހg���ߏAbT�ɴ�JS�
���/�	��`���W��Xi���$���� Q����ׇ�C�}��lM�e?sř��5����7ϭYe�`�H$%mt�����.���Gtt��"[+��$��q���l=�o�6�Fo���Փ��^���Z�I�0>���������l
��x����d����.���)Y�ڳ�fҵ�
��QroH�L5��o�u����*72����r�R�P�H�}�����`,Ӭr�G�o,0e<��Tm:ab	�L2�J��w_zkL~AN%t���mIogM|���2@H��#o�́�рT��.�a�����0��r2������l�r��I�����,dmydn̜�&Zq��K��j���4��2�!���6���?�^{���<�ܡ%�zō��G��`� �/������2Y���<��3�\`��fF(0$O?E�+���f<R�Ky���C/�h�K"?
쿟ػ�o�l��n�pb�mP���}u�ʅ�չ���8vi�dE����7�z{�R�8����(�����8�dȥʭ���[���c�T�#�t�+�׺�� �'Dy.��f��b�$4t���!9��
��uYp��Ng�4�L�����{��4�I���E�BjU�λ.F���)��r{�)��i��~� ��!q�y�7AI��8��=(d$�%�ȟ NP�L�us����z��/��i ��{�K���z����<L�l㸈�jp�,���i̪�@�������2��2��H?��2����Q�K�~7��&�qU�t}�a�H5�ۤ�p�z|���q��n�H��]h��GX�gJ�P}�B^ˇ�ƣt\e�TC��E�dE��?[f�2�*-�N �4��߱�Ʀ�9P�|����ō�o��ĵ�N�*�&~M�5��ܗvF��J]ɛi��e+�7d-}no�a%,�b��4?�R�1��mRHO�Ŗ�G3��Ƣ����%�5�nA�z'�[�b| �>\��hw���읭P�lc\��|G�%o����w½�L�)�EB�|5��xF1#����Y���Z�C �[�ѫk�iT�'_&�#���<�'Qq[ �thtۍ��i�t����qȔ�B���,:��r�<�����ۍ��3Y���棫������ݟ�{}���Q%?.�xbؿLm���w����G~E~n�;����+L��j�֍��V_2~~�:FsT��͊3гk�O�݁D�F�9��n��p�G�c)�Ш@�6"C_ۏ'.�D��M� ���-�����)������#���C��� �߃P��<֎�DY鶚��E�f��fr�r��f5v�����7L��B��s��L*d�*�B����xw4rJkt_�dUl�c��:Z�²�6y��`~��(3^'���`����Vw:pvK��֬XtB��-���O��MK�dN��h�N�P���T���[J_d���0�c���(���E��]nD豇�Z��b��)��a����?�!J˳>Ea.�d�n'pu���R+sO^'��P5�K8�p���g����D͒i_�ཝ�	�Z0�嫹P���"<���+ism�o�ͯ���iJL�*�[	
���Iw�J*	֔�U��谵����>c���p�t��<Qޟ����,�`����<��MƵ�u�['y+ $�y�?@9����~�V_X�uR~���]u��z�40��@G/�x����%mw�M1��y�������闘*�+,�#JNE��[V�ַ:�-s�\�_���n���8T����4��	"Z����x���o�:�ফ�iob�ƚ����~�̿�S�������]*D�B Q�2�{hr�6,"��q�&��*ۜ�Â�j�Eô�p<G�iZZ�j=�*��		��$����hU}D�����X�`�vz�:ƾ5Z��G;�ɾI����Yg�MGY�M���Ԧ+��E��ɹ����J�4�b&DdP�O׏@V�a� }��dY0mA�MS�R_.��.]
Cp�Aݎ�7�~?)Ict�T�w�@��.:��0aw�> �'֕(���Ӓ��ӿH�X� z�[���Bc����^WCM���da���B�c�Ͱ6DG ��g.��`�I�+�9��q�%��ܧ���@�aܔr0c&��Q��lt�\8�]��d������E~���P�/���$U�-��0����L�E���GE	&0�V�n�^v�R*�8`��G���hؠ)�4��
����=�d�*�̙�iͯ�<�����("ѷG1�r�]���ʺ�}ޠ���X����	���7��\��de�]Ri;y40,�;�=F�u'4��x�@�߷���Dp�.��T��*e�-�
�8��]��D*9�	���o��%nrfD��3vv%3��Ky� �E~������2v��zڳ�ga�H�w95u/�N�1�9�"PՆ�����z�G��'���[Ӑ뗐1��Θh�ȳ��"�܏<gD�����,w8]E��z6ˑo���Rc+(�;뭛#�^��L����hp��qP ��]G�����&&��|w����%]b���le�ϡ�ZcJw�QU%��V3�f��~�@8˻�O��G[�;�b�9o�˘VU� �-Zԇ���e�{?:-;9%O����e8͞��w����Q;� i�R[�#����������,���\Ui�lf}mm�Nd�k�g�t�f{���	��-�%����Q�!߃�X�#���X<����
�1x�9e#�;�9��=ذ�j,ͅ��I�G#Z�����\��%F�A��ڰ䃳��ei[��m���L|*o�0lS{�[����>f`�Kl.�z�g�.�@V[h��-����o�3����?ӨO�+6�CʾfK��6ņ�/L(�9l&�# @Ƭ�����NG&_���Rͫ��wI�����Eh����U�U-~�lG[>��WOO����[5-�������K�V싧=]���TڙCK<U�T���
�� �f���Z�v3ǚS���{�?������`�s�\�T4�=JԀ�icr}����:\1�>h;�9q��^HW��"�:`ީ;]��kC�)Z�1X����#�#'-E��)@�t���H��;����/Du�x�z6�Uzj$�ǁ����ѫqD��1"�����]R�M�ׄ�6a�qB
��+��U�i���η�	�Y�^�� ��]-�a���QB��	t@��Ld���K�.T5�
��(UL�����D�t-����.�`LD%�W�{cr��&���;�sR���r��F�n��R�qM��kRA�79�v_�;��c�9}c�L���ӼA&��j�����gh�
"��ٟ��˽�\N*�����9!_��Y����Nv"I�u�����,gl��G���b"\	��XbH���P��8O�Mķ�ʶE��ɧ�EMy�Br�I���D9M�G �;�?i�k`=��(φƘ�R��$׬���
@��a��j]��q�L9��V/�F�w��]KD,������a�B�n���&w)# ��mQ��Ot���N�fq���LBʑDB�z�ϩVda�?s&�GTu>6p���Yڱ��#]��9����E�ʙ�GIm��q[,S,��'�Y}��h��
J�lۆ2���C���>	wuo���踍������L����nhaP"��j��T����hH� Q��ݘ�2�$� ��+.H���'R��w����0䆦�auK�%�K���p�˕,�apK/
�mv	�u4~�e9��vں�Uv����!!�	Ʈ�43�!�"x����Z�4��ev'T >Z�!���p��E�*���h�?���nz�x:�?Ʒ�~9��{`^�N:;���{>t=�|����Z[���e�a-��bs�D��O���ή1�h�[���;�i ƾ{�Ƅ �C�i^�Gx>�����=<:9G�������h���zo��Ar܆����f-`빷+@v�B�vM����s> d$yy�}�[C�R�>�YJ��\@`-T���u��ۧ�~p�	ׯ�v�Fu�H��E�}B>-�i����ͺ���������;;3׊DRwU[�n���[>1��b�l���|҈΀���s)#�w�����^?J�%_!��®���������춬���IsH�7.^� l(>!/���Q1�F���W/yu��Xa m
�hI�pN��(P5ݕw���|F�˔�q"���9�&��?5s�1�1H��un5Zs_�nk��.���oa���X=$�	�G�3��n���ˍ�'��X4aq^:����̫_eg[G\�7�"J�̖��.���Q��b��^��(��7����vԊ67|L�䉠��	ɑ;�e}4���Pf�{~H�.@}Z��U��d{Q�/>n��rة��a�s$���W���.�::��c�&1ސ�P:�ayh	�Q��y����M�f��[5��
�����_6�z�=Y����/�<���7Y%����^��G�1A�ȹ J�V�l���"���9�ڐm|YH�;��9�IUޟQ_���@��d9�N�mm(���ݴE��
��w9�5|���թY�>�;J~�vhL��?�_�l�Y'�F��d�8l�Z\�5E�h��Ϛ�}Fv�~¼�E;�QD"/JхHL9�n�Cm��b�;�ܮ�ˣ�#��;�lg�hL��F'��PK���h9sd���o���G�؛+(B�����! Zk��挡@��IĘ�C�=!��bW@"��TG��s(���Sa�g�� ᜷go��k�U���f�3��d8����M=����I����zӀs
�ص~<u�)�E<㣷CÍ��<�,��QL��]��$�������H�x�*��j3}?�iI�H��F!��>�!i����\�U��^s'���c%;#lI��8[#ĤU�^��e�i(�À�ӱH��t�q�E�{�Ŏ�z�'v���|DZs�r����cR�1�ȴ���xHG������|�ç��v��j'���R����Y������.��#ĹL�zy�no
�ݞ�<��V�4�k�"�,ADv�)��0oL���ys��-9_��E:C���Ĕu�/��c czC��eO���{�St�9�lf�ݤ_�P:Z*_��:��Y�/yɽ�&w=j>O;��@	��1�I��3ݲ��U��{c� ��nhئ�h��:P��67��"�Z�D��?�=�q��7q&T�A�V�?J����qs�haQ���2�	r&,�?��$����paǔ�W���kk
�Kq�-X�P���-�d`������{�P�a�z�୲WLJ.]ی�X'ڶ��zq��	qx�>��;�
����$n�uv�#⩠IW�+��!� �e�*S���%���]��?�� ���--��ڃ�G�J���fk�������9�������A��G���V-��Ӏv����ށ7(�\R��,���`�@=V#���`�ċ��+bc���WX!��&J����;����Z!�P��K������ҪoJB����_�`@�|�p�UZ�Ap��E�O�I�Gh�vTc�z��\4��Gwh��l�OiS��{�.0��o���/�0�D��4�@��NNXe�/-�O���@�lj|t�|�ά7���a�������/�fզ�cU����t	�3d��o�iTI�����V`�\]F�4T�7*z��	�θ��۬��h��8/`�sX�������p� ����9‗������5��۟��z���h���Տ�2��f�(�7�O�!��V|EQ5�s��*ef�	�����@H�C�ѡ�^s����5˭�>_gX�Ϥw�F��N�`E_	��s[����J�¢��:��l0�`�1QzG�`X]a��5������S�gG�W ��M�C�(�O.xD#Z@s$���� AbP�&̫\R�������O
N^V�t��
�H	�Ð���0P��*ɒ��I���մ��n��¦�mO���s ���#��b����v��?Cv	/��րA���n�I���1�}^�Rʩ��Ќ������y�Pk�: ��v��%<�۲e�U�����k���K幝ղ������Bв���&�K��C���������+����~c-���g���bG�����i��ÀU�dN ��I�
�= s�q�e�X��mܜ|���Y���.h��X߈����^X���WQ��xcz��c���J�����������W�u��(�& ʸ��2#6-V�����[�~��~�L���Tݝ�s��' ��%q;��C\�s&�<О4���D�4�tt
�9�:��v��b�k��c�Dv��~�8�_��͏�_��d�g��`][�u��a�d]*�˂�9i5#�6Z#+��xS��2�} ��1���F�\s���ʎ��BD3�F�]h瀠^>�*$"��1Y� �>}姄��`�L~Ɩ"wn�2:`
��wb��j@�������H����D×�A$d�	_���h!�"�%�.��E�i\���̒�.��2�䧅�����?"7ʠ�g�T�Fzi�MS��o�܇�]ig2����"��;���Bh�tC��)����V�������\
�O
Cc�H����(��m����Q�B��F���6<�d�(�
"�%C1k9E��y!����;Ox�U��E~|�ka
�Y����Ė��*�)�7'��n�>�l� ��|�ܹ��ئ I}��mB\��%���S���I��2_yg���Q�61/E���̫
��P,��BO4�}�.��~��6�X���(j�^�"��&�/��2;i��z]�B��XF>��)�ҡ�\��'S~��ڟÜѶ���IO�H=�[u���N��:�9�&9������%����Az�Ӧ!����Uo[�_f��2����Y��2�,�����$\ffw+u:����R��4Xa2