��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv #�@���i�\��n�A+A�d;[���WHn��.�w�;63�L���ݷ��K`
P�W��Eh^�X8��S��d:����/�{� �'J�|Ǒ�]��ځ9�)�vM���{�9Cj����>�b8���eN�ɜ�u��F ü���g��=����I�ʒ����N�4�~�+N�b������wAٛ<���8摟'~zZYA�6,H�ΰl\ �	@�9�Fq�=���!���M?a3�XU��w�߱�R�H�E��4D�S��1��Bb#�:���"������fT��G7Xk����?���5|6`%�S�$�(�}�������P���%��XfºO��a=ܒ�eDnrs�.���ۜ��m���'�JS����Ԥ�A:�����qh���,i*��X�]�N�X����;�* ���2+��v�gj�L��U���^T6��,��	�����^c�N�'�e�W��8��N�ɼ��(���!��U���`G��弦��1uBu��tN���>�;��d����	!���/���ru�0��#>C������V�U1O2/��/!5 Ǿ5�İ�#��ҏU��R��V��QSFܝ^�ʯK�Ġ��Ugs�8:S}# �KA%1��w��R��q}f,+�Q��M6�7l��+�ѫ����܆V�(��CIPcz{��[���}�L�x��ô���t���äI5(Hb�g)����贿B]@,[�d�5�'V�9�ƊJO��<��M��կ�}���^Jv��K��E'�*I������Ӓb�q*��P����wM���F�ѻ��r�j�������EQ�аAA�{Ҙ&ZË�mYe$j�I�~W�BOΠ�)���}4&�%nu�(݊kA]�G{������g!�~�L�.?(^-�YP%QL��N|�LI�F+�¶{O̔O"��w�?�:}SW@0kQYMS'�2���}rނs$�������E�R���ǿ�Ǚ7��ܼ��v��q��@m�6(sdMw���)|���_����O����zqü���$��eׯ�9�Swp�ՆԻ�SV�D����Eޠ�����1����A[~�@�`���Y�o4q��J��e��%�+��|.l���+n|.����
>�����m3c/�����	������I�L/�}Uz;���r�-u��[�,�Yc�A��E��\�>�J�<c	j5�>� V̭9��M��t�G���@�).ɯ���-H��o3Q`_>k(�g����C�6����Q^��HT/�>(���܉4K꟯��/��/��н}�u��@�2��v])���}1���t�L�TX/P����.s�Ͽ!܌�Q�F*�B�88������n�2x���s��I��<F��=�Vz�p�[萭O��<a�A��|��<l���y�(;�;���!FW�����O��r�y�.�Ԇ��#嗚w.�ZK? �+��r�ȽX�X��M�	�X�ƣ�<��i�w^�jۨ�me��R�y�,Z6�B@ɁB�����,bHg�U�`�[�g��wl��� E�߈�ݷ�Q���RPoH�3�.���x��t3K��P��A�S-��{��ާ�#n�+�@��<r��*���CU74���'�d!����r��f��Hؙߧg�FKu��m&+Ts.t>�唯W\��[�XMfI�X��#����c��j&}���u����Z;�@|��4S��˔C\���A�(��̈́�Kk�'+����!�;J�m��B��?�a�?�f��t��E����>Cb�&�m!~�Ѝe�||b����ȇ��d��sp�����"���Y:����TZq�ٶ.�h7/!x�A��`J��Ǹ�J#�V uel�xy"
�Û��d6ܺx���poi�Y3�ڟ����J�K�Ve�UP&I�����:�ZYX~�`,�)�l2C��"��Ȟ3���K�0L�t��9�*�<qs�����~Vß	|g���>���uX�:�#\��&D?7�q��ӟl�揨���L���U)e��w�2���ߊ�^��I�.sz�hj���]�X-�%4,��1L�v�)
X&��K�؆s*�ߙ�i�z��� O�=��f��r��s����Z������rW��'+�qV<!Q���E��`BѴٯ��ʣz3&�0>�l���0?������H���Vi�	a^JR�dK0MH�.�5�t�d��#�_����r����a�4�ʯ���j��:Zٲ Q'Q��&L6&_uq�(ԆK��#��z���1^[��#�n���?��o���lч�8�}c�wo�%�Y�J�yQI�`ʲ1	���3�k�\yC�����=�=9�>F�g:$�}��*�ґ�%�ґvE�h�̮n��E;0	����$�R}?,K�~���&�ۓ�A�l�Ξ�*����u6J����4sN��Qd��7�jy[V���@��Ѩn�}4#`Ӓcцַ~7�n��G�	�*���@�X(��F�#�h3�.v�!�lw�V�ڎ�v��ҜE^����)���`�|~��x��,�)߆�|sP�.�w�Y�f�}�����04��{�~��Q�@6��"H�)���F��	[�N�>���0�ߠ$|=Ɔ|�� 9�2���7{Zo�!�u����dw�����u�$&��S&���.���g&"��N,�':�)�ϞwC�Q���.��1Nd����f�Q��_��2R3ch6(=׈�U���P�9�|A7�G��<�ȳ�j���E˒�Y��~A�܄�Qy��)l��:�[>��ʁ9�!��3khQLp>������l ��]�ڮ�A�~Ϩ �ix:�2�$6g��T2�H��a�i9a��
���kL�/�A&)���;H�o�9�o��AtY���t�O*�b�
`����\ze��B[��%	���7���s�E8�ER�_�� g�q��K6�����_�k��ɵ�`*�<�b�%_C �^4Ib����`NF
�Z|w�v1ϏQ�����o}p��	��a���� D�S&�?�x��nYLmg#�@�΄Θ)t�� ��5p�6��ș�^Q	���L��8�o��,[{\TZ�W�ծ�Tcho�Y�����C����U�0��ly��S�[�%m�(�a�,��A3Xx!��Ʀ%��i�1�OaK��U�R�s�W���l���ҿ����[d�EƼ�"S6�}�<o�8�����$�Cc`?+j|��D���� U���B��������M3��a��$��
��7o�@�z�:F���1Q�����QŸ":��k'�|FU�*��H� �� ó�BO��T�<$�<R�H,�]�#3L�#h�o��x��|�Σ�#W�hɠ�F.������K��k�S��>@
� 3JW�YW��\����CA^�m�=P�(�����5uN�g�9��f�����!iNLLX ���0<�=�|"-�Y\=bׅ.G���j�&a����{�e��H�����(��`���pl�8�_5����_�Zl��ᵏ�&�[��`׵��CUZNё@�E���{��Dɤ�a�k��v
Ŏk;1v`�Z��Հ��4�[+VS\��[�;�S^���Í�p����#9�:]�Hq��n$FJ�U�����̈6���t�Ȼ�5�~ţh����R����ؼd@��l9�R.4�$��KCP��lݗAS��=�� ��,�zs+a@<�yj����v_�n��K���
��xԂ=锘)4��ϝ0{�6�'�������`��ͫ�f�����J>�Z�!�T�zn�������r���)xDl�z�p?��r�[(��2I��-H���<�6%�'�AΤg��'�o� N� ک���L��9�J���zhU�v~`�a����������������~��U)�`7ƛk�Z�� �-��������n���\�~��&8����b���ނ��=۸ܮ0��XNt�%�lݽN��*0�w�����t����c��|�T�<��kS���joj��DI;!['��:�̿Pgp*BX�0v��c��p��|��-�oE�f5g�Q�e��HE>�C6%��땴k۰},ND�49j��탒D���N=��b�_ye��K=1�U�i���0�V���KYeO�aIiC��X�}ݪ��ʚ7��y&����S��((��Y����P�}������I9���|�G&Tw&�O�S)N�,mf:��(������[��'�'����1X[�S��?�)�m`�W;{+ڔ���;}���bD{����q����u�;���4?F�`lw�h0�U�Sǩ	�FcfQo���X1��X�Ľ�ue�#�	N�N&a)�|�壩�?����*{
['֍��=f�SOC�Y���c7)�7#$c��F��я!��$MK�ڣe�~������h����&:�wՈ�6*�'���4C�~MhЭ�b�_���d�&-��tL���l7�Z1���<�:;ᴸ}Źj̤�:��^N�Ĩ="-�}	����SеAnq�⩖��S5�/t�c��*3{�n��Thl$A'�u]������Z@SdZ�5��F���3h��8�����õ?w�8��v��a��E�b1~��U%�n�]����Z��l�-�(�i��A����/qkЋ���_)9����'U�@]�W����Na@��V�Xc^b�'\`��Q�Ȟ�w��oJ��%���?慵�k�fF�kbb��6�u��� *��㝯��Rv�:]�\����4	�����4Yx�V����j�/"�����{i:�9@��C~�#�[]�FH�@^� YX��%
w��d���I��"�{����^@/k�|Gw�8ʑ���8o�pļ���;<��=��TҼ�	�./��I3��J�p\���ٔylE����= [��m���H����`g41.��Ы�Ͳ��-��_�#䏢������4���&��M$~;u@�2�~�ʲ���~���4�f[��E����ƍ���>�Z����4"Y���s�����__���7 M"�#�\���ȱ�0 }ٚ�3m8pL��=h��WKv�&%WB���\WBk�U��=��ӭ�QBf���ޣ7iT��<(��U;a��i�.t:��$ 0&]7<M���;ws�>��y&4��xa� I��\���:��^�#(� �o�B��*T}m�ѷZ?��6y��Ƭ�����H`�2���g5TtB�F��;����ݰ�������r��,�"�YH�����ĕ	�3�*J*�!���߰=+L�W�Dҡ%��i��妓\q{�핱�߮��#�.%{DDB T�F��@qC�=�^+��Tl� �� r�&h"/�t�M��ڵ�%;�ve��f���w"պ�p��J�3�"�e�E	8T�M+�p����n�2��L�ѫغH^HI&m��Z�T���*���֣pfѨ�L�����V�r�~�$�0������6���@��n��t���~�1�!��z��xq�Y	�����@�g��m�kv��V�O�-�DQV����\���oq�K�o"�4,���2�q7��q�M�_�-���X��>��k����d	���6�7~����o�;-i�!���Eԍ�
jh)t�@魴���4]L`EY�%L�`/؏1�t�D��>��һ��/H#�/��;��h�Z"}:�Z',��)���+�S�+�G��8� Gأ��L3�Bu*�p4��ϠG����r�G|���*5N�4���p
?���Dy���;��uۡ�O� Цn�;�L�������$�RS�ۈ��=����{��	�b;}�p��G��y�$�UU�]�ĉo��J	d�����q�@�3������jʢl9[��J�����w�uR�x�v�SWT�u���J����W�AA�k\&
��wîJr�cڡip��+,�T{)��� ը����V �� Bר ���e>��l%�*���>v�Ƹm�t��Pm(��An���O]�	#���*�ǜU<���`a��tSGs�w�a�k aTO���/p�u��m��� 3.�Wҭ��iQ��7dP�5GG>Φ&p���!kd�$@�\���(js�)�����\}��������U^��.��ּF!qv�X��m�t�����¸����>�4�N�)��K�\�1j� 7�$��8�i��bkN��i��SY�/w��� [�l�P�Qj�����r�#B�F�����(贖�k?�:w6�&��nΨ}CG�A����w�ޢ���qꄽ�u�$�G7���'�栵r.��ߏ@"��ť/6����P����Ӣ���t���V�fA��![)'B�s�#�T��*{a�&���z>���(("8mc�#��J(p���`5g�ݰ-�*hm��Z�t�V4\dD�cF y�!�O�Æ���{��ʏ�D$�����N��!�E��N�[=mPz�3��Je�ݸ���Iu@����zc@��|�J���xU���iu��<Y��G�w|�����zX�z=I	���lv��@�@�2�ۙu��"0,2��+	�$L���F)��.���6tg`o@u�a�b�~ :��P: ����e��fzE�� 8���r��1�Z� }��׆�kb_��u�sv�h\��J�PQZ7S�V����f�ؠO�x�g�����3�%>BF���q�aWl	�'Ɇ�=��a�Z�N�����j�Ë���`����/��������A�L��(�J��3��n���+�$�P;ĩ��s��qo�^�X��&� �+P���9"w�⹈]��_}��]\p�@?P$S=���O�iLՂ��A��\�+���%l��
xwQ�R�F]蕡�����&a	�wp�����������^X�S1���������A���5�XFYR�B�ɏ�F���B�-�w�A�~<�}o�۰�p�� /6�iĄy��C�+�<�� �c)B\����b��)^ɟ>6hH{Z�h����Q�Џ�2O@�� ���CS_ѝ?M��fp��+������/,��>J�q�FB�#� ����j�_�,�����2�A+�V��D/����K�8e�ۏ:��l�Q9�O?�m`٭x�ĉ@&n�-����L[eP9�\��	��m��l�1�&#�[���[t�F�L��uK+�^���`�1�qT��8G�v�&ĵ�"opQ���٘T%�=F̂3��'L�6H�����l�C0�oJ�&1���-L�_d[m5����G�=M�1h�?��!�j!�2�5�?ۭ�"�HL���,Q��*/9�I���5����^!13��ͿK0�.��q3|�ʜ(=��*�L�T�/�`�:��T�����٫�|�]0\q�خ%<V������n_�f�1�/o�^CSEDp�v���`�Ru��.�Y s����[j%:&}ȶ��*�6Y��nON<oyr�$M���ە�N%O5��
!	�Q��8����&(#î�d��ݺ@L�F�Nl���	�.�bp�ѥ�qc����V�W��i- ��z��I�3;�|����W�ƸƁ�j��p��n�5 %�O�zie#H�7������������GU�E��K}�]�T�NX ����8ׇ*E����,ՁT1�>,S
&D�'��6x�j..x?�n1R�Y���!)E>:�w�uBO	@ɦ�]��47��p�{}���?i}NYn�����2�����?�4y������g�~{���O��!F"O\�-��n��ix�u�7ʉ���h���M��x���SM���g�k���d�}�R���xJ�h9�s/Q��﷣U�H&Q��NærS��X*�n��۞��WR�8Hx��l����R�65�2�tṪ��/���]aN�u��X��f���c��}�j�h�ǀ{��"J�WQ�n�x����o�X���<�abuV�Ip��<�bg��Vs�����#��%(��ݨ0�_�e�r����67���b�z @��2t�ޚ.e��V�޶�pyqkkj��(�r�U�z�.��rJ�t����g9f��jsL,s�3<~C�R�T �m%Hv#O�1s�L,�����r8c�;V��,
6������SR���� �ѯ��oߋb�)�t����Wo/�&:B{ԗ����ɠD�(
��c��|C�r�#��|����gH���M�(�I��3�dq��Ԅ�������i���P�-=�ᐙ�8���?I�V#�VP���顱�
�ã�> �c7�]���x͠�-%7�!�d�zj(�{�%娤�Β�ە�?�R�ϐcצ*"
z����F�)Ǜ�c�u����h���a�4@/c%;�i3\n�4������x�!�ـ�?E�A�}�6��BvI��9+�2���f�5��L����v���f����+��5;�N�_��1�x�O�
��`��"��q2-L�t��	�L�����Z���C���d���U�fR�����'ݦ�ؤX7c�^{D�0���tv����뱞J�(ɆXejE�K�����h�W�L�3�ڂx���>敄�ᩐ�[˃������G�L���)�k�,K3�=�撾�.�B�y��2��d-����@�0�p�5h�c����(VGib��4G��tC�����C"�T���N�y}�ޣ��9�rA,���? ��Ol���w�%%��s1�_�oeZ��ҷ;%�;�#��A�p��Ko�&�%Enܯ<�i�W�����Ϛ�����V}X��<�8�[hVj%g��~���e3�a�8���N��cI�7��ȾR�� n��D��Ȟ&H"Qrd�.2�fp��͜����0�m?���A�f�|n�(�VT�#D1h�nPgߎ��\�v]r��	�c�cr�R���[<��k?RI�M�|���Wd;;}f�R���g���σ����L565a�+�j��y/I��#Mݬ��J��ʢ�X�tk��oV�LIjHN6M)Z�Oۋ)~�[Y�\?2���(H���D����� {�����}ȯ��&��D������рJz�i+$�J�ҝb�?�~��*�;7�o����n�UP�9� �������-N,Ҿs^	2]*��@�GY	�8ꍙ��b�"��N*�%p�P���V�.���Z�9��O�}KG"Ȳ���ߙ9��I�G�ӭ̦儧L�� ��ܰ�{�R�̛us�^U�UB8��)�θ��s����t��{���LB	v$%d����x_V'��ܙ#�����2��6Hj�f{t�RD>�ko�Z2W�B�N��]*G���yR�I/�ǖxN�_��C*�?�`�3t���0$e��N�|N9$B�i��g��J��~XO�zEx�w�z	�J:�f���G ��� {��'Œ s��f��*4�̣��#������U���06��J]n&�ܠ�Ώ�~D%��۠�4��ji����Te�fޯ*ش�&J�2�+��O����a%��ߺП�KH{�8��Z�·>
_U�f�{�?�Ǣ���h�����͓5lܕ�4�UƔ� ���}X'Z:�W�3(!�l'66��C��@��c$}��y��Q��߶�zuߝ�M��=q%�g�S�=U�ӛ^եbB�挛Q��������n/\v��������VQv#�Ԡ���'&�Ϲ�icG��d��q-�X�o	�������=�Ն�X,����/�~*.y�����N�OI�o�E	��x�2��O�k�����7݋�����?�k�ۛJ�f[�EO���[��Q�oH�iy~�I�K���u�n�7��#tS:�]�����ɯ���O�,�)Mv�$����p\�Q��3Rx�s5:]��P9�X�;e���)�\�)p���K�N�C8^�k��/��ۻ��6��A�r��<�%��|��^ޥAa�"��lM��mrq��M��O���8G����ļ���h>0����4BG��u��9�Y�Nr�;!��P��kB���i>���erL��C��^jw!g#@�ꏦ&�u�Ґ�12�RW7�:'��f�u]��S�( �ë.]Iu���l�rc�����C/�v{[8�b����=�_]y%1,�=}9(��~_k����c��r�2פN��Rk�!�U%FK�;����0h�5ÿ;��B��DZ�8��� �斪9&,x��U��
�}�]/��(�aZ�����������P�/�ӓ����Kfbjd˧�y&R#��3��>�cR���+JTK3�3�-޹���2�H#vg�R�W�K�@9�}�^;LgXv剑��?7VXW_�#uk"�$���> wU�]�K��F�cJ$me� D�A"_���9nF�G�|h��#���F5P�p����~(i��QMv?Lx4�0{�=Ȑ�����A]�Ax��O)-]��קX�A�j����vn�OKS�L������4x�J���ƈ� Ԗ�$U>#!�Ճ�.d%�>|{�����G�u3�·��������9lgt�eIg��{M�Q<m��a�W�v{oȥq5{k��Ř�冢�.Io�O!��!�m׾�"�v|���iq��g����}���, ��%�ΐ�6PW�|�(�
; �{�J$����v�@�h�n�;��&W����^��U���p�S��%r�ؒ(���4��-I	X�ťe�<��k�͈ޯ���$UZ�ύ���:�VG� �l�(Y���Gp\�P>�4W���U�A�KxyȏJ0��&�����\f3�|z�-1�y�e��;��sHF(��=:�U���>E��cu���r��5nڛI&��2��-B����sʦ�)/^K�u���C��7�v(�=�p؋��|%�t�Y%s���)����G�G~����E�/�#��YG�_�C	юj�kO���.ri��o��c���ԆC��J�% q����pS��*�W8�|���S��0S���X�~���K(8�q�O9O �p>�Z45�!2R���2m�Z�F�E��z�я���u&�Q�J�≛J�`�O�������s��W����i�;c�!�]ϭ-�Q�;���>�Gz�H�.:.Q�ۈ��;�X�J��r[#��AM���"��Ho�%]����S�g�� s]p^�⨅gIQ����?���l2e���|�!GKٴ{g�`"pu�n�����v{l��zL?���I�̒��[{Ȝ��w��^qu�;�	1�a��T��E����	�o��}�kX�4>��ݾe+ ?�V��F��vS�#I����U�SƦQя{B����2�Ѵ��@�
s���0��)��ЁL��I� O��b���"U������8�"�o������Q轶�:n�C�� �s���Q��癯cZ�,eM������|�z��'���5��6f��]o$��y���=+�i|�jH���{49�W���毲����DP�c��8��,����wk�T�;݊�ɵ;�A���A��ޑt��zZt��n��A1�8:����T�|�d�O�,]pWrTGSz�b��7@��pW�ˋ]9*d��]�%AeaF�Ϸ��SUe�����0���̃Q'��R�!��ZWXa\�����Ā���]+�>�cA��5�L�D�hL!����6uӕ?~�_�L,4��=����(S���"Zf��3/��}<m<@����[���%�-�M��/�R�
JB]3��ӯ0�DX/�T����x0�|/��V��ZV����DS�/�+�kPhc��̭K� İ��"2��n�a<ۡ]�fU6FD�ew���E�& r��6�S�ߖ���4@(��s�tP����#��à�#r�`�K-)e�X9��2(�w"@��|$R������`�\��������g��Ƒ���qm<�Wu,�G�$�0���j��Dڕ�MUً
/@�[�`�-�`��bR���%^(
~	BQo\W]ot�]K>8FiP��FC���p�`I3Vv��ϝ�����&�@w�=r�����������؂0	��ON݀9�+ �O������O*Q�s���{�6�+Ĥ_#��ӻ�;�`lp�=��X#�zXi���V{j[f����,s��i�%�%�P$Ы�s���i}��� ��%�L�ІD���>]]��g��N�
]�i�{j��Pd4!U������M*	��i*X�#��8]��PŁw��&?O3����W<�5�F�7���A&��‾0��@���w�����t�7�-�o��!�Bt����^6&���M�k�-�#H���W��Ӗ�~P0Ur�a[��n��5@��Q���Z5�"������[_�����3�$�!���k@97.D����*���E���YsiL�'�ϲ����)͜Y�63��,,��8R��,;�2���OJÇ8��'Ã�F����/�x|nv/�$3��ϩM9pE��="a�rc^n�/	
�ߔY��4�.k{�3��RR��k2��*qOͿ�����aI���.�(xN�����h�����j�WPG��MU�
��������9�bKs�kcL��x���;��ZF������/M�B��YŰ��V�F_�=풬丸���C �t��D�D5�!��K�U�Z&��1��	y�G�|�ϐd5E(�^���.�&��K*	r�'/�P�(�6&�@��g�H�����+X����Z5q����{P����f����g��;�t\|ymL�"M�����U4� ��L����k����SLiqC�e嬜Q6C�a�	����eZ�Z�j5�J��^�n#%R�w_S�}1Cg5���C�1�Dw
�B�ұީ�V��fdJA�ڷ/.����5YOD�����Z�<p��ŭX�IY��� ⓋW�	�8�;�O��y7�2���������ą2�n5��A�c�I���B�U�⽱,}��J3��v���[&�S�\���%������Y�8�hc��G���ne�0��ȥ1MV~��q�pv��.�O�(���D�a���]?�"h�����FU/̥\Jw�9�LR{�)bw�B��q�ݐS`�����5�hAM�6[i�?o��߆�V�#��6d9�}�O�v���t# ����	���^'h�ld�
�‶����ܲ|�[�C�;�c��3�$��r�}+�J�Hk*�uÄa㪬2�IظuG1��Ik��,gɶ�(a�y�� !l�薀[`;��&�@ـFg������$(�Nc5�Z7H.�(�K�A�<g��9�J����$\�������OI�P����b:����d,�<[|�D��<���γH�Mw����Ho���j?A�|ޢ(���fC�*F�0���Lr��J�R7_����.���S�ۇL�@��f�E�K͎���訤CƢ$��A�jB�M%��g�j�lk*W(\W
�,]��F:����Y�7C.l�7���:��S���>M�����q���C����\�YP��:NvM�Xcff�Htv�]�*p@|�UzM�%�<�@�@�����z�bd�$��l ��-�o�f����{(�.#�\v��ޫ���@������4.����Lk��b�ZΈ��S��^�#��g7�DÄ���ϱ���Aq����D�� P@;�vph(;L�Q��F��j�ys�06�����ѣG����+.�O�5����N�͈Ľ?-���0�e\�>B�Ȁl��N�ײ$�d��4��5`b�(M���)�`1[J���#�q�H�~�N#�ThFK
�-���yBu_���ˌ�į���Z������a`��o(������]�~,sN�&G�{!��k{��ȋ7F��O73��u-�/���T��nJO��Z���^.^s5�6g�)}��,8���S�?<\L�CC��௻���k���K���b�LU`�a	���Z;`VA�ߊq�[%At?�,�ǃ3w�9z(@zi����CZ$�a�_�w{N	J�e�����<�`������?�vh�K��%fP����%[(�aT�������Wn���v�or�eU}a(3�wi�nJ�;���c��saЭS"�D��<eI�K+ke��w ����
p��W/Q �a�[���qNVL����t�4QźL
�|���X��v?�{n*�����#�}(֥ה
���*1�$�Ƥ��e�ASu�O�U]�Mֳ\���͐G0Ҷ��2�&9�K�1kd��'�۽i��r�Z��g�J�3�S�W�T"c~�T�
e�֤����yg��KBG�
�F�I�m�ȵ�� ZD�>'@���C?V�&g�H��&��9�_�>��������l���K�3Uae<�1RZF*�>���3�zF�@צ��  ���>�
�%�7'w��s�U#V����q��Ҷ���-;׾<����@����S����q���CZs�趰��nhc�8�3Nt���oX�`���K�f~/8���K'��� ȧ'�g����IC�b:��H/���g-�2�k�P�݄�c�����_��(Y�&|��ŕf󧨲�o�>�u5�An$��rÖ]m�7��l���c%���{�����d} ���$�l�M8X����H���"���S6������)�c����nrI��$Rj�������ͻÛF�j�5&�%/'���Z?S���^��F4�@N�ci�giT8x�~�9���R���UX����\d`��-K�v�+_��x�F�_f��.����C�9�U�s7$8����"�N���,2~H�x(�/"���1�W�K�[-��.'�ĺ�O�g~��
?e6p&���^1@L))���%7�]�"�rLH-���A �&04����a���	����5@�"���9�$ҕ�15)���*�x����;�i�=@o/a�M���s���a�E����@�"��IG�������E�y� Hf������GT�M۬��ɰd������AX��~��>�4��9'���p�����0�����Bf�3 *�/%�>a��ю+e6`V9��[��1Pu��"��1���'��aP	�-��om�6���R24:��z��qx3�s�d�D3E�����-�X�_m���l�j����Sa����VMS�ը��BĶ�>��
�[ݯok�z�:��*6!I����7{D@���yq�_t��/���$���ao��.����T#���6j�Gg��VDE�/�w-��t�O�s���2�6l^Z�"F�a�>�I�@ۋ\:�G���H7�U���N����ӓ��$����@bh���d�a��Z1��l ���l�A���Lܺ5dT�����l_t��䫡Vtd���B����	V�}�!z�����_�
y5��}��D����E���\�o�Jb-꭭�LY[��i��\���a��3��ȅI 0��d��HL}�58��>���b��TYJ�FL��^���zU�O}��>�����N���X�\�Yl�V��rhga���ܯ��1%�-���X�@���իH	��/lg2*M_K���r%_o��Q����C	7Oex��7	�Y=���=:P�isL$l��%-�nVj�
�G<Qh4��{	�����>�£�eOw\}x�%&W�Ӵ;duUe�9�{�Aw�
�����R�"��m>�'��]T����� �$�W���}�����V,1ru�W��2/��n�}P<;Zt5�K���ӎ�Gg:*E~.'fr�"!l��b;�c?<B�Q��A��d�^��hPjܼ���t}Ygvmd[�m[�l� �����2� ��	#��s�pA%����T�F�����Z��YB;TRm�.�༻؂/�K\v��8�M4�����e��IAy�}�jǱM뗱ϗ9$Hkc"HLsi����M�U���7J��,Ç��;�#�%�l�*��5�ʄ�������̃,�}�h��,8��!��X�Z�mW�b��oM$�P=����"��S˼�G���IK0�[�t�\8ڴ�*�G�W������kc8�S$�ӝ�"x0偆����3��L�O�D2�����?���q-/U��x �2��&L��$�ڊ�*z�튮�):kx�F� )�+r�cp��ow� TXHķN]�Σ��y*,��2a��u�T-�R�+
i���z�8������M*��H�2���u�|a^�����zO��4ۏ�s���d_LdftC5S���́~�9Й-����A}����\��i��[�<Rk�ÍَA�@�/��:��2r'�t?՜%�}�����-��t�֭�j�C���q��Izm_�(Yh{�� �N1�z�� :���[8ti�b�^ø���d�<��� �o�I��?��0E�%�y	Y����}�OV��WV��CZ��5�n�����}�!�D�[��^����)
��L§�������j~��d����D_]{��P|���5���n���}�,)<�C#us��{_��<k�1��C}�x�����![֎O�%���%O�l<Bs����VD�򸛊'{ȧoV������F�(8m�c�p�Z����M52�x�F��y��V"�� \�.�]��T.	��X�=1��C˿�)����E0����fc#-,�A��/^�eԲ�&lPLؙ���M�z��LH}_�l#�+z�����9�����S��Z��5r)�d?�
k/�
��G�����s���[��v�S�4�N��6��UN_+0��=$$�N�/ݸ�؅�� ,�3lžc��*� �C��)�8W�p��$t#r�a���"�ߣU*2ð�6:��=X����Q6�<N:''iT�T
��H2}qY���9D\Q��t���ł/2�Д*� t����*G�A�%G��F���gp���W
���� 6�2�����NZW����v _�P���o"�q�Yn�a�t�Y��Lxm��z�O��>pHٜ��_�z���V�$�ѽܕ�{ ��T������V-�4$�Q�u��o��ZE�]�V�Ȏ�.J�8�DIm��w�+�~6!�U�ׄp������#�۔���}�.2Af]�W�K��!� �tJ�T�Tp��0��n����Y����9�j��Ҩ���O�W���|_T��-o�o��7�No��&>[�}�߼ah'���th���� ��Vr�T�>���:��njlxǙ?|���5iΖ�VD��G5L,�]�[���+a>��������,ƕ�1�ȡ����H<�'�L��.�ҥ��-���S�j�Eu��Zj��{dI����R]�,�d�W�����Xm1$��ߓ:8b��m�������r�@5�~St����z��A)���a>0'�}~�AI3�kd�c�9�F��ٺ�M-zcU #~1^��u����JD��� :9U;�tA�I
V�
0��;2��Af��Z]�;/l�aa��)� x�B�_��c�N�W����@zԜ��\tj�9>y���R"R�BKQ �A��z>M�
1��v��Z��D������E}Ɔje�1��X�]9c�\��$���il�4�߿�;0vO�wrEN@��d�Sf��*[�1�=�)��t��l-���˄ɺd��Nta���yIg�ع\�=�x�A��|e�
�9I|R��| w(����.��MJIT��|�*�=�R�g����zɩfE���s�Xܵ�JbS��%-�u��&x��4��.̩���fD�[ Ab׹�B�m�-��q�^�2�-g��9<:��/���1��=>��yH#_��M�>�!IquF��׏�S �B4VOo6��'�pܣk��l�3MX	uq��'1�����z���3�01�ͤ�Ψ����4�ƶ���m�e���ټ�FU�.W[>��=�(����$5@��ie���i���u9p��"+���܆����jIξ��+�:�̬�j��F{G�d��0L�=�����I�~d���2�8'���	�la��L����ìâ��nb�\�3�R��oݞ���S��[�/����V�(�������<R�'�b���+������KU�-���'���aE���س��FBM_���լ�0�Z����Q@�%m�8+#�Y&H�zz�/_�?vxUs٪����ý]5�ǭc�Ȍyc�a�8��v�|��ԡ���b���vι��u���/�1����`���jzQ��x�&|���8v�;מ����L�Ԝ��~F��cB����:����J6p���ŗ�	��^�n���¸���R��w�e��s���5hwV��j=&`�Oa���O8�`�8$���y��N����Cj�����߁f���]��_������u�[t߈���Z.c}x����?ĥ5���2�����?��^���
��#ƪϮ�B%�d��=f�k�Y]�k�L���i��@#g�b���A�JaD��s��q�e$�� �J����99��ޏ`ůѪ 5�jͬi�8�l������U~��U���e5���nH�ꑠ�g�>��zˢ �&yԗ��)�SwXC��%����Gp[1��	)#�q$����1O�W�Nk��+3O�6^-D����&�Óg!�[����Q�L��t[��c��k5?��k@�I��,�<3�7�8C'����q����Jy��d�џ9~�m|�o�L��Ӗ�g��s������U�L|O]�u�����kl��c���?��,D_�ZF��XɁ7W��P���.ȠYE�Y�A��Ҹm�i�@
)�/d�I��*���A���`�P���>@yʰƏ���������T���΁'BrZ4#�D/�_K<+��{����=�^T̶�-B�� �-�vw?{ƷZ��Һm\����j��$�?�ˡ�޺HВ��Z{�����ZJDw	L�) �����?�~/�d�R�!V:�*��Q="����}�@��Z�%J+������gt�D
�c0[�9m��}��aAI2zJ���hZ{ml@�v[R+�Uw'N/`1��et�'E��R�o4�k��#�p�H�섲��3�)�n�HO�A�_���3�]�au�	_ፗ�"\7��#���7��1� ���D`���C>�M�|�w�ޖZ͆p�2�%�q�0���hF�����v0$
��0S ���,+�o�רMg�1}�,
ȷ��~���Rz.6���~Z��=<���m�dn�Wʣ3��O<"P���ka����y��1�y�Ԁ�z�_�~���EʩBt��jڟ���읇�*�,5;����h��a)�-ލ�����r��B��w���B���f�1\��������"ʟl��B' E|'��)I+�_�����e:���7N�A�`g]�܋h{���$���l��ਇ���qՏuq�X/��b���:�c���pӠS�D`\ST^š��.��AJ���3c��}bT�ƴtz��q���p��֏`����\;S�78�q@�cvd��w7h���C��~j���ںsKw><wdۣ��cl`�ydr~�������$����B�7Y>�,^��Dc���
4i�@����E��m���T���&�[���Jy�������Ǆl/r(�
PS0��ERؿ�H�gM��� |,.yD�k"{���ydk>LQ�2�\�f �a#�=��z
���QÝ�<q�Q�T�y��o?��NU���(�&/.orh����2��Q*T�t@���!0�`7/���,A���މx:��.1�����)hv�B�ko�?���M,HN8��v��[l�-T�3�s����ZWE��A�F�I�k�j�P&�d��q �.O��H;@�~oz����=u�s!/��:���Z<} ��*u)����4�Hih��㲲�WT���\��o����Id/�I��g���b�v���:ߞVI��å=;�6��GKJ\��U������V́oI���x[
�%]I#ӑ}�yo������9͗������ayG�#Ъ^n�C&*�>S����r�>��Ŕ���%���
���D�~>��LF%�Y���d����h��A817mhG��^�bȝ�[N,��
�b�H_�E��.\�Oˬ��ƒ�����~�P=���@���u�(��*e�W���+b����a?_��_h�I���=)�C'��.Lp�.����|���N'���G��I�{#{���Y�aߑ�>٩E��b)5t�ge���6�L)Dd�R]�|�c�e�M4���T�`P}���O�l@-�l��$�
��V륈��I�R>�$��27�8��S����Av�Ln)[w���CD��`Vl�iA<p=�ٕ/K��`�nX0��T��g���Ga�H���pגK`�#������)��n���w�V=>ϕ�Z��!�o�bd경90a��o����z�׉1���c}E�]��E��w� �c�Lw��7�� B�xUt��.R�P-�_�K`w̓�>�h7O�+#������џ6�<^7l�O݉'|30r�_;��ڗ�1>-�d�=����B}������&����R@�:�-�v*�?�.�z��s�<?� ��`YϮ����>��Cy��9�k��^)�S�M4�YG�|q�[�����i�����N��yH�'�ld����uG W&����qG���K�+��Z�g\l�����2��_4#غ{��	�M��V�б�ކ����s�ǉ��E�_|���e؝�'ƻ�����'��^��ޭ�Z및&ٲ��g-y���:7�$�P$@o��$���K2�z���n����~"C3p�5'���}
Pxx'�Xa��)�-��	���4�{a�qW�"Ԃ2�e�s�^59y8ҕb��j$��*ĭ�j�o�}����FK0r�ܰV��!W0diçSIu�+��-�R	�9����2���ӓ.����vt"�d�!�f[�|I�^=��]Qp��Y�� �E��mb�|[c� 	ץ$����FG�ˀ��P�.�/�>搛lݩc��{�!����ZH�2��4��!=�;� ��5,k��o�H���\\̷�ˌG��=܄d���_��Z8`�j��/@��7m�>z
9��w#1��`,�!l���X0��*��){%
� �#�"j�2�����f}}�a���1>��-�\�I���-��(�+^o�f����G)b@���k�=�&t/H}I���*���g��k�l��B��:/��R�t������l��V	�����B��I��K-z/�cP�YOjL���կ@��7���,%b}4⏩N�����ٌ�.�7�H�����<�f~����c���I��l�g�~RL6^�g�%L꛱�ϨR�	��BopR���-:���j7��1��-$M�>��sR��D"��~����b��c��N�kxY,ԯ5֬�v�b��u��O:������A�f����k���1�eK��&��3Q.'@�ϕ�$�F��"e���S�JGx�LhI.� ��Q�~��R9�SA���Q"T�Yع�Fpi��+J��31N�m�
��:Coq;���fks�|�pV)��G �~�i���	K|�_Og��D�Ln�^1�%�\8(�pG�g	�ux�/g٠��OF��.�j�m�P���U��a�Y�߁~�����|g^%'nKԣ�a@]ח�np	D��N������8����uŸk��W�(,�,��9fN�(Ld&���w��L�Z�%�hӶ6��{5� 9ڏ��5�d3�b�u&W�Z�z�G���z�T-㞟GF�9Ru�F�(�=�\f�v~��3G
圦�2�t"](וq���?'u���8�c�) g�D��]FR'���<�n��J��ۨ������+4�ֵZX��T�U�Q)�;�Z�p:�K��5J:����(O)�i�Dㄶ<�Ք�7��o�qZ�4�wBcf��\�� HOlП�=q�3m�-��Z��Z�����l�\4��B���Ӟo�#
�Y�l�.ױ��¼��6�yş'��9��Бc��^��Z���E��B)$'M���O/)�>�'�1���?�ˌ5ۄҲ���'��R��@"rO����Pa.��ѽ�Y���W�ލ�9@"#!ig�"��ni׎XO,�:_z�Ҫs���-���BK~��>���pY*�j.��Ho9���G{zj{�I��0��orz�N�C� �-�]��k��t;��L�l"�(�$>Z�� ��[�Wԍ�M���y��6⭊T�"�K�Ǉ����D�"ŦOD��������j��;�2�~I^�.��[��Djf�v��!�?�����̄ ��ӊJY��W��Ҙ��H�)ob�PP�8Z��1E66K�<M�3����b]�ϪuH�`e`.�[��[���H){�q���ϫ����r�����2��ĕJB�Go�� �b�%єa��do�*,�^��)L:�]8�����nM�8����AJ�`����Z��WgX�~?V��B@.���3�{���w����wΰ7<k7kt