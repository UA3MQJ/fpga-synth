��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�������V�B����(�1��~��Ԩ�.W�������`�G��}t�G�!d�\L�q�'ʋݟfe�m����;���܏����w%>*�o��Hi^oˏ��WA٫���Cټ\$^1@��Xj��`dP���
ma~���H�JN�y��th�ڈ�|�*���'{E��; c�R��l� е��|og�*.�n��Z� �qg�=]G���ȣ������TF#M��u�l�s�,1%o�]�M��qH��N��ʽ���dN�z�T-
8%A=u����6 ^�xqF����z'���%�A���q�
Gk}h3,��[��u� GL>����C����+R���PG6:��\���;,c������KU�#P�m��J_�����/�)JŬ��2����N�ԍw���j�Hh��t�g�G�"<�	�}�s�uB��A�K�-�ͅL�e���I��l��B�&�`qf�w;Z�/<G�&ݎtt��� ,z�Ǉ��=r���v^�*�^^�<�Y�G�}��^�BW��W��H(���C��o���K*^���b6lfQ��}���<��T����������(��)���bO��s�䠢'�
�/�sy�H[���PO��Hn�]��̉(�՛�Ux�`�8�C/��)�}�͆��L`����_D[�k��n��g
�C��*�ρ�)g�E�Iq�j�����*?�vV��Ѩ�|�hA<q�N0w:!D��͚��ۘ���tM)��v�!Y��Q��(XK���\�K��8u�O�xs�)� w%�*������$��d��JSi�+)&�
ow�}�e'��!(�N�_)��?	���z9�m\@�z�h���053�}�I<1,�E5z��E�ӄH|�#�R4�6e�У�8uaӏfu2����˗߻���ZO�(oޛ��N;@z�<���-;f�oZ,�1�VC�t�"ZJ�e7��|�O��@�n��̺�<�q�!��I�Vs�����
�u����st��Ѧ�ɸ*f0�����q0��ĀP"9-�J�u`0]����V.E?~&E�M6�J9(_�R)�yy�w��ЌFN��f93���E{�'X��ɭ�4,���{/�9��uwaSZ��A[7:��uM=�*N^H�cF�ۆ�^��㩾Fz�x�3%��/R�?P�)��c����J.91�N��2,Ty�g_F�C:��6]p�8ttsֱQ���B���z��X���ۍ���7��B���t��O7�wY��i1��ח�ho=�ƌ@��CIWʽ��� �רژ__���T��kؤwT/�?�
/��Q$����5�K�kdT�����&�Fu�2dTX�Q㊶��;�a��B�v5��������+�<;'���W'���	o'������71��x�����1V634���0#����}�{9qv�D�yI�T�x
ę�Mpd"��˒g��@�Ii�YY�y�*4��9B�=�?���P��Ը���0�TG(�ʜ�]��V໰���\&�ʗ���"p6z��
ub��:7��tһ#��>��Cl*��a4�_��]��J9��b>�9�4��w�ޜ�lǕ`(���D\���,��T'T 
o!'����9�+����x��p�N�*%�r�个�U֋�l���T3>`�Gr�Ǹx�ZE��B��:H��gx��YZ�d��	ȘR��l���i���F���䳥۔�����2l,ʥ��0kf�8��\�m��kM{�����L3=?n��zW�1�(I\�|Bj4TnM�L�'�����ɡgِ�kG;�wA���9�/�	�HAA��ݗE���� ��qX��*�s�p߁�,��WpΝ´\����ebx�`#�e��Ɣ�E���9�ypO}Wt���|�I]�"ѿ��M_�#�;F�}�@P�#��q�
mt2���\�J�؎?r�G)}*��z��X7 �o5K������	�B������ �m�փh+t�u��;i�8���V���k!� �����FѸ|-X��٬I`���u��������ƥ�4B3���'|ӷ�c�E�������p��,yhe;�&L�sp��@���Un*���0�׊��cd˅ �7/�noxQ_C��n�Ύ/��]�M�Xn���V	Z�T!f�#j,�b�ؗ��$��Ec ��G�J�.���yp
[t���
o�>Nmd;�!�op�����17��>�u���z�����D��GQ9�}�0�}����Q�$p��w�r릱[*:OG�P`�Zp�|Ew'�ʷ���H�m�]O ^-a*�F��J���?8�v#a��K4��k#u%}�c��d��}��n�}8�H��)�����Ymq,����=��P�HoL9 ��Bt%��6���b�\3;]y�Ďd�i�+��B�J��Eȣ�$`��ӹޔ_�MTKٻA��*��X�� g���O��ܪ�ڸ�Et��<�^Bn+$SZ0"Œ�;�u�8�#Ym�Ɋ��hj`0�/�ڡm��g����m���i��G��g���?� ���ː��p<AE��WN���բA*;zW���9�I��&���	PـW`-��f�u�<��S�M7�X�ݒ�Cޜ�~��>�+8�nF^��m���8�>��2jN+�Z�Cp��>���ϯ/Y�UT++h�S��)Mk���5�=���bʲT�1]�p �� �̧�ZO�*W{�xz>�w�vŲ�d\=T�\#gL���u�~�m�����&�����WiD��� !�3�m�� ���(��e3>&Bbt���Q�Ҭ�nAX�(*����<�?��6|ŧ���C���L�3��>����'\���M��7	A��r�`X�@r]R������_�xJ]A�L��Z:�|NzWI��)O��wja)m;8�ĳ�����8-tn������!�ɀ~��TtX"���YQ�ǟ�K�m���Z����$E�i%��c�P�������;E�7�H7�Q�\�c	��IU@.��eg%�~��\(�m�d���v.�1�v	>%EB.g��~�ˑ0fE`ki���� ��5Fe�f�7��� ����Կ�f�gė�o����%,iDlmH ���E2��N�5:�K�q�K��THz�j98���E*�ʭF;�&�,�@�9�l�V�a2�QjWK���! �nW��z�k��UT�A������F�vm�db{99�84CD�)g��	c���tTY;�W���3���`���+S�I=8(u�R�>��o�c�����3�Ca�Rn�oms�*�o��#��YK�M��n����@g.&�>�˘��I"����L�~�=T��@���L��P�̘~E�TK3�S0b��mZ��?$V���3Ӈ�AK5o��(Q�U~��&�k�5��_v�ɑ��FP"���Po���c�|��ȦR!T8<`� ��s z��D+�Z���$�"*�L4m��O���S�	�A���dfS�k�c��=�TaF�Əa�.�u��9K��g%F�/F[��E�s�	K��?M�#۷�ƶ�2��$�q��PV�HEa5%�w�6�*dg���D��C��c������u���O0������v��=�Ǽ>��r�H,"
7�[?[��U��4^]O���D�BLT�	.`|:�Q��2�:���rB���	�F�y���nM�:�
���gRp��Arʸ�����(`�J�ʗ�"��r����D�C��<[�
@#�A�����7AG�ĲW��0�x��qu��nՈ�r�z�
�A�������3l�q�������P��.@U>):���!�푌}�L|���p݊&�a>
�A�j�5L>�x�`Ggޯ7�� ���m_�~C�A捙g�y��&>N�� �|X���2
��`BVe@r���?����6n��3@��qe�G�ٗ�%��jqό��9�-�4 7n�*�:iD��{�w>0u:��<r�zS7�v��+�n�����Yk�a�0�����Յ���S��񣪓�Ȭk�:،)+�	���(�L�]HHL ��K�����ƀO;��E(�*o����W�[��bWK� �X����9c�=q_�=��=>22`��aK�Jb43b.�:��jC\l�&w8������3P>��+�����E~7�g�͡9���h����2�<�1�<�M���>hF>Z�tb�|�pLk��@|l����0����d���٫�X@ԒIO�O<�w$��i�k?��Jo���uP�-��$h��6�Oav�P6�\M���Qf@��Fa^(��O�Uz�ٹ�\Z֘�tX��`w��:t�,���ND���dX%�Of$�!�|se5X~�z�*ە �_�=;]Wy!�l=���$�Զ:�P�k,���0�TKOIn�}:Y�ͻ���胐�Rݠ^�8��0�]�;#�V���\�x��P�C ��ę%����IxBv��7��t!T��([�r�����I/z�u[=���j�@��_����f���9�����{��m� -�%����EhI���K�}�鈞6������9L�JD���!m��1=,�.j�QK5�)�ӫ�ʸ7��@�����Gg��I���$S��$�=0��z��$�	�K��&Ï�p��w<vnc��joF�w:�ը��.���6T�w�	z ����u��_��$�5�s*���YY*K��?��C�����q�=�xZj���Ŭe�h7��5������O~���9;���!�;��	c�o�4
��Zk���/m�`���g�"o�����X驥�3�����7�Nm[�Tj#�8ce���
uˇ;��x�T!3��]�H�8t�������~1��.B-���-���`r�v%��/����|<d���W��lN���D�a{������a�G7�tC��z���OG��Ƥw7xF�ϗl.�� ��/B��PׂXD8{�l۲�}���\$.�X����;�7_b�%��"<��=�"�Q�9_�Z��Je��bS�W�7V�"��)�B���%��|R�H��[�j��5FUv5B�Ed�TXֳұ�AX�W���i	~����U��}]��&�nH�A��)lHE������û�Uӛ�u����W���x��U��4�
O؇jh�ؙV7f���ަ�`��R;�Ld�o�� ������6��W$�a�Mp!���/B�F�Q�f�ve�*�*�}M%A���Yyk��k>�JR=��f�kP��Д��^?U�����+������.g��D��HH��J���^��)�G�1u�|,�1`[.��S�&M��:��/�"K�]�7N>!E�D���c��4��B�����j[2(�����4�Y�"I��S�2�{�0��4��c;w�/~D��u� �&^5�bmd�֞?��ni8���N��U�@���@�ي�~�����e}C�Pr�_��>��qV +"q��T��0�{���1i���k�"J�4Q���j��6���ѓC��Wj��ui*�������nԈ��9�'��tAF��|V���F�X"Oi��I�\�Kp�����pw�L�S�
��Ґy�
��s"����%���s�L�]F�:��eK_�<0F{fn|9��½�e����W�2(��&Ub��_�`����jb�(�Nz���w)~(�`������<B�-��h����|�77��x}#4Y�'�@O�-�	��̓,�6���F5<B��
��J9�N$����6s�zΜ3 �3%J�1����ֵ�}$��kȽ�\�E�N�T-1�ΣT3��J�9�����Z$ӓD0�ޑ��/�bor��7.�Z�)��V�E �nʗߟQ��˴:��EtUw��d��DV��+E��v�8D�^`fM,�����
��z�$VJ�������n���!t��s�g�[�U�6ml�^�����+�\,�?�5��Ϧ�&*��J3����*G)��ي{�fFr>�N������ڏ�}��ް ��r�9)s��^+��2P#�o%�2�D���p{$���h�����O���[<���ń]Ȣe����W����Bx=X�0��W��UP��5~3�az0�ho�)=���@��?<�a$�N}�m;�k5.<L6T�?�4 �ޙ�`�P\hA�r� ŗ/=f�e_���<� ~�k�/���X�5���?uG���q�d�&F�尺dH_-����Ԙ+�Ij�W�W5�1=J_WoO�I��g(��
xP�,/
՟���%Y:�:�/2M,x�f����kQ�z��,�w#-�1,F�yW��#g$�j�/r��)�e�U���=��>I�Gj,V'�3�
�7%�- �t��[�:ާ֪�������U~v�a�F�!U�5JC@Y�vuT"�^����V��b�)�Z���y��)fۭ��+������QC�ȥ�.]���B�[��g�M�b~p��2�'zRd
BH��0��8`����5ItD��@|d)�p;z���۹A������u��Oy��ǡ;b�X$b�-t�?�1 i��]��&s4�B�@h��_�'O�{a>�O����s�h�.���ى�%Fm���|�r�D�c���]��9xMְ�s��qQ�-`�K�s�;��e��]Tp�R�X�e����v�wj"F�������*]��d2�S�kDĊ(�2��+!��ǹ��O�I۱��l�#�I%T�3'X�,VPS ���c�K�p��,1���b�{��f��.L�c�i�,���؁����(����5��^�!�[�{�t��t��)�)��V�Q�35��|��ʦ6�E���I�5�2��b
{Uu��N��Z{b/�X��qYE[� l_�<����y�<�J"�|VK{6èo�3A3��+wh�{/�"�1x(}�=yÞ0pSh���J����4� *�=����G�����@������	��f=~MaY]�-�S�|���*�蝂�x��D��+g�㭉lFJhj�����)����S�$>e��;���Z�()Z7��0�+�c����^#w�_��x���E�4���[��2�i��P��4_��%��Q�pt��*� �T�� ��p���n�?#H�8{�ǔcN����m_���w�.ed�b]Д~�f\8ͺ*3�RE����e���f �cEɾ��p/9Dછ���$]�����.��#��bP��yQu�7���`%JZ���&<�0 ׵i'0
�π�:���˂+�x`Y�16IӮ��E��(��u2N{R�s%��iA�M�W���y>;���>�ď�N��5ۛ�1N�J�Ғ{V��Pd�7�G�3!�ՃS�si��M�&I��J����������SD���t�� R�~܎"���Q%�	���X��ᇋ!3>��w��	Ʈ�b�X�����b����e�zM�����!b̆�3�5l#� v�C}�J�@G�e�K���>A����ȏa'���Bni~�����2���	u�Em� ��<n9�:�^��&x�=�Ȟ"��*�/�U�bv$�n���<	'�u6$t�Xg�UAؙQxb�
)���>�����3��qW���Z������;��`5�λ��/9���I�*�g� Z�o�f	>G��.�N�x5���K������:b����`���ʐ	�;|Q�ߎ�=�oj�C�e������_�x];�8�ó ,�Y�a ��$��(��gM!o�����BOe��~�7��]'?��ͦB����#q�iV���z����jJs�h�}L�!���{̸�K��n'i��!�~m˭�q�Zj7�5�>C�ϣ>L�Ht?�NV*L%}�"����|������F��򪎂�'������^�ò��	��B<X+��+2}�D�젱-՘�q�l�8$|�{��<`�%��8�O�]�'Ц8���$��]�֋��8����?ȃ�.\z��!K{�EiJh"X��_�-��a���{�C$��G1�[��*�(�Rq�U���8�à_P�^��BlJ/ӂ�� ��r�1�J�������=�R4E�;?�z���X�Z������
�1^�~u8�˲x?Ԁ�-�,Zt����M��dFg��h!-[�	�1�zթa,��?��D��n�-= �@Ⳟ��D�?�@b�
��Z�^�B�%�ք�m�9��dk��E��} s`�{�	F\�(��̣����~i8ЫNK����M��9+����b��Y?��%��fc���4�L	�g5�˻����U�x�2ˍ����4-6�q㞒��������7R�sk�����SN�]��%f����b�ܚ�lXn��|� �{�@���h@*� Sl�������'53���pA4����֘ON0ۧ�^�{�������g Ȧl���.ZK��S�G\�K��^}��Q�sJ"�Y�e�ok�."c���v�O\xL	[������ �x��ty�DuG
+��	y?�����SWX��/�^����@�,�Ȫ����q�]I��0%�(*&��ɔ��~�PI�y~�Iӄ��Ī�\p`� P<n2~#7:c_�H���7������.o�r��J�����v�J�n���O�c�|�n� �Vs��<�l;�.؎g�fQ���C�?o��U^�m,�|$��"�US�-��:�4dr$�lg���S�)�D��U��~��-;^h�b�)��(�g�kAt�
r�X��d7g��ÿ�`�ճD6kK+�.��>�j�(����\��X1�re��̠2;��-���g�54a�-�M��kn�!���_�Ѳ6�\�o�J���]#;y�Y�5�9y�:���e��@�oL_��=C����e�o����72y��t�̫�	�`���A�e�f�Jxk���N�8�k���w���|a,�X0L�(o=,BТ��Q��z�L�!1-�����B��ݮi��G��3B�%����앒�9P��j��ҷ�7�ɨ�����B�N�%�!7��®;	�@��a!N�L���Q%?�>���� �!,�C���
�����X"P ��K�@8��7.�R��["|��4��Pz�}�ؤ'>�
��+z|&���>��<�p\��G.��`��Z>�J���'�I޵s���@\�f�he���� �X�]ݠ�Bl�������� ��(����")�y%?՛��K�^�3�<��!q�o���F��Uh1iQ��:�/�ŭ� sS9��w�h���pQ�9��RsR�Z�'����|�@�8����հ���-L�c|$�懺Z���:�S�q!���J�����-El�s�a���7�����Be��EI��[�`����i����Z����(U���[`��ʌY1Y'g����i���a�X2��x��8����y�G�R�?A&�J0�h0�!���˔�ߛ�(����B��L�ɍDH�2 �B�z�p�g_3qvB�`4�nnub�E~-[�S�ʙ�l�J���%t�	�{�}dio��g�E�76�-";����i��o�P�nH�I��We֪w������^@R�F;����������`2�!�ݗ�-��~��ܢ$2�/a"2��1-G�`6����Dx-֔xY���6J���ҽ���7&�wzj�D��Z2?���X
;�b��	,^jZ��#�@��oBC�I.T�D%�2�<?��G�u�9@ �C���\���(^���i.}�Ÿ�"ʮ�OE�*D�b��k�c�?+�PF^�����y+��"�j;��3h ��H=O�!�B$mQ�����b��K���{˿43�k���)
F���S��k��A��]^�A88��D�U��I��]�1`';��т�-�hs�d����vǦ�P*�Xy"��2��CЈ:��CǢݠ�-�����+ M�8�s�&�ĈM�r�*��A���ȧ	U��J��4���;���2!a�9EĠ�>Z�hV����a!B��FY{����˾�4�)Z���/�c?p��E��* �(xJ5]�*��J�|�_�ٸ��?:n+�P�b��{��ivH�Y�1�½����R���A�u�4ݼ��(�"<E�2��#m��G����m�/ӓ�A�ʧa�KD5�o�>��]<�Kb��O�Ř�g�-y�Z�<{O�4�3�� _�[0�4)w狢յ�u-/���w����� Y��uM�:P�(V�4yWy�M8��*�e��2p�]��R/��<�)b�DkcYzY�'��hI�U#Y
 P	FO��۠�z+w�{u6s��j��7���%)�r�
�W������31�aH׳pE�,�����=��	Kn��J��Ш)�x+Ș�ҡ*u��ꩻ�0L�4�՘d|Eo�L�gY\���o�yi�kŎl[��W|h�;�a�} �����"�#cT-�L<Z3r�m��!��|!���;iS?$=�x{�d�3?'S(ߣ`��%R��M�����(�b�S�Z�N]���9���
˥s��'���:bʦ��o�Jl��Y U`��!A4�m�GlxU���1hIpH��ҧyX��R�L��F��˯�����yXLYFB��=�%ۋ�<���R�l]��1U̦	���?��;�ŝɎBM{���3���߭�fÌŃ�W��MLh^����H�Q�a�֬ɴ�y�z���O��⥻d��I7���Ag4�x�q�TA��#������mEX��NY p�\�]�(�P�5Fo{w䢜�IY�ׁ��n�r�|��
��r˒���*�5� �zU`c�oO�� �Q��m��ߡo�ǜa�� ���B����L�. �d���Zt�����h�y�R1�˥[=y�����I�D�cc�\�El��"�o�1��[B��a$��0ZE�q�G�]����N�~67Y/'����:ֱNPq��w��yD�wƬ�\��0,�"
1�`�fMu|q�/a�S)ctz�8Wx��)͖�1VP����#���r�'8�ċ���~#��8�B����1�'֘�xA��c��f�z e�*e�t��PA�I����x�KZꕿ]�� �J�X�e���~N�` ����j}���!�n��Q�*�tl�I��B�[aM��G��9Y�tE�umx`<��o����2��Fi��@���7H'	�W,�p�]�j�㔊�&	��Pr�����_ok���N�G��"��H5Sԫ���KL���c��nzaH�&����1Z�<�Z��fl3�?��>N5N���a���1G���8�.�U�t�<�:�]�`�>r��PW ����2f��ŚDV�GZ]���,O$6eK�[5(�mrT�ܱ��|�}B8_�	���H_��H\����̊�QN��� T��wr�3w��