��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc��3@���;��̵*T���që �|c\
��`P��o]L̛�鿕Z[<eLl˭�W?�;���Xo����^����Z�<�F�g\CT���/4�Ǎ�@�����(�Lx)�EF}��N�QÑ�*�����Zf�ϏJV�E������V�M>؆1"��0}��{�ƽ�`G�%[�,s���>�ӹ*����ںA��j�'j��''$���F�Sy�,�v��i^ٜ��/f���.�n���WG_�kQ
-,�.UI��ۉ;��Y��ULCͷ�,lY{
��B���<�����N�CĖ�Y���3r�����M�Y����1���{0FN�_(s䌶8�M�QtB����̱��GNZX������-�7��&qt�:�I*W�=�'md6��p0�F4��/����P�C0*4vF2���,���ub-A0�����A���M����&�4�����Nz��g/��Vס�%:I+<����s��w���5;qV�fȔ��ȟS��w�D�ױ��M���D�k�E ��K�E>�8Y9땪�8˃�t�Ϋq`̀h�9��8:�A��V(�YX$�Oɬ��ء���~�/�
���r)�Pe:�����Q�@G5|D����԰��jQ|�7B/��
�8"��3���P�^�:�'(U`�����
7�;8�M��[{��l�nG{�f(",a�W�A{�L�vv@�9�Yk��R�[�`�qbu~���ٜ	@"�sZ��4�X�1�k카�WT Mȡ?a5%��ݞ��[�4ח�\r~bW�Z���R��"��y���"S]��FA�4t%���n�H��o����8�(U����.�2\D�ۺT�oRՇ����U6�7����z������9��ke#�r�T.�\@�b�B�����H�<�d�oa`����Y�:0X�K�Y�x�T	p�!;.�T�g���b�K�W�G��C�5IibHsC(J
~|��O�
������v4�r���W~di2`-�=M?xM�!��m���X87`'2Dx0"���~%��Z9�c�!�}dfxe�>9�#0ܡ�p��&�@�$���I�W�A�&�L�j j�3��Y�`[�G
����w��`S��g#!z�Hw���'L��&6ׄ���B�s`$.W6+		�6��g�X�+��qy�`�{�|���CS����j@�7q��Iʼ|~)��G
 �y ID/!]6����8z�x7)���RO���O��گ��
����J!�a�8eȼ��:s�OQ�ɏ��\�,ў�G��FgE�;3^^��R2[�����I�\a�p���l�:&F����&�
���Kqf\/V
�w�sa! �P��V����e�uMYH(!c����ڣZ��c"��~�H��Vy�&>���仆|��?F����������R١J̹�2@~�.�qX����kZ�Q��tY���f�i^w����*�[���1����"ԋ��Dp�[2��Q�c�HrZ?d����$A㙓T����Ҏ1�r" 9;��w�z�H*��Il�7�kS�A!��g}iÞ����,۠�E ��E)����{��qh�*�ZT��-�)_�u�9u��$�R��*����d�)�@��T��n_�� �7����K���X�S�;u������I{�xJ��W���5�r�񷆿�O��A˳�{�Ƅ����(�M����@fb�}��!V� s�d���/H�w�5V+.�?/( ��r�����~T �!�c��c��N�e4��X��|C!Xw����1��B����b���ZLZH#�:�3�G�t�����k��W�O������Ni7�׏���\P#8puA��{u��a߲'��8�fS�q�Rh�ʚ��w��+�=���PbTI�ZU8�'*�e������F7��ɻ��d��J�I�ɢxj�~�"0]ʇ\��N��z�[����v��$g��Lg|]��Ò��fe��h���|w��%�|p)���W5�0T�Mq-���_TX<w���-�s�"���@e%~(!���砂
箔�I(���mr�+��I($ɫ6��.c%d�~��=K��s�Ʌ���yi�ξ{J|>l�'j��^ey�����dS?%��EG�8U�R)3�X?���!��>7���2�9�W�����pq���pʐ����зg/�EF_�Z���_ϫŬ��e��Tt_w�Gpx�7� �p�}�6��v�v�}¨�d��3����'+~RWU0�'�pR���O��8xM�M��<Bǚ���J�GA��v�и��۝�\`�~�Gq���Mb2��u>6�hs�.l/M��`(���R
��苙�W�%Q���S�$���؏��ϋ��N���c�䪏6xG�qã�����O��۔�~�1�м���񓛮�w1���[��LtH�H�}���LKo˦g��ʄ��/m�x�u��9�Vc�q}U	�����ذ�dd�7���L�O��bȿZ�\�I[�6���s���3�̕�zX�9�;�$3���<]��f����m��>��L�ɝaZ����@��ʷ&��ʰ2xb�$}Ũ �f��0戍ǃ6��$��g^U��&��n���!�Nˑ�
9�N�/�T�}��4K̹���}t8��a�s���%�&�e�Ӿ_�S�?l��Y�;���榪�gp9�%�G&�#O<��<������N�<k��vF���D6��{���C~���)�,;%��PmJ;҄����� E6o����b��23�z*��dFjQb��^ۑ�m�$ks�ǥ�ۮ�ъ��'_,[9��uH�{�o	b�WT2cY${�#%fc.Mk�p�g������h�7@T.�[(����a4)�)��y����U"+��0�1I��`��ސ��=��;�Ǒ��+&fN� |0u:F|�}��3�U�o����i�j4�R������b>Z���ī�a�f���q"��^ezvT�i�C|4�xE���ܚ�