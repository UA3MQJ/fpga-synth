��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^(Q�`QԤѥ$Us�fӓu�CQ��rƙ��t��uī3�m���j_Kn���&Yp"8��_�X���qS�������~x
o�{��0v1�N�^��uv�N�S���@:gW�����ם?��S Q� �8^�������?L3��j�+��ڎ����Y#�3��X��\.�#Y.DӪ��8�WkOo���?dJ+E|!�3z�E��t��z�s�ۛR��#O?�{DJ�l EJߐ-'���3����F{L��d�� �;[Hn��jy�"�E���si�嵙u�}M����G�㩠_o�߁�2�Ŝ�<v��e��A��K�'Xs�D�5+�����K��2���ͫL>_��N�D��Rzʛ���G@H_�Y�����"8.�R��-�L���]��)x\�`�(sp�L���(�G�;��
���DW��g/��+�=�͛�h����l��&�n�ܨ���ɠL���m�8<g�@A2v4����8�z$�}���@Y��n5a#�8���	����9k|>�~���TW�6k�4�����[�C8@jSy[R��|Vg�/��>�t5X�ūe5g�ֵ����U��Hķ+ð�Px� ~�3�.�/��I��-x����_����`�(���f�Ԋ�'���C�o���3�r#Q����8�������Q��sp+U�^ə�;5bNG���e�5����Y�9w�d���6����������8�S����R���fa���=��sP��i�?�?Oq��ոo�M��;�����u,!8+���Y<�*��m5��[���K��pҞ��g���C�q#��S�A5��eq���0X���MO�>��s[.���!� �BA݁�ғ^��*�	i�!u��5A�p3��ΗPX���A� �������8�yu�1�F����D��b���G.;�-�J`�M��l�1�>z�R �0����(���<�9�08���b�u
�Ց�φ��zpx��}���"2�1H�k_�:G�ͩ�>���4m�:���-U��8�%֐��$'	H����/�Z��C$�0�V���A��0^���k��OUﳅ���oD���Q�,�S�������{/Bu`��MR�'J��D��g`P��U�N��s
qy��<�OSOf�f��#̂�`M����UOC-��o`ZC+zS-����Q���ا�pCO��H�Ά>/?���'n�����~��~_���P~U
C�?V�I�t��a/I��b��A�!�؅�HpG�]@�@��d,N���*�<���L�̻y&���i��֮���ڒ�vbtvI[�XM�ǟ��}۹i���Z#�,2�q�}q���u5~�;�n��Y�u1,H��^M��z�*��5���$���;9���M
��4QO�/�V٦�g�����_ .h�q�������8��{9��n����?�'�p�*�܋�Y���97"#�b���<�r�H������z:�yek?��50��D��X��J �c��&/x��3���,l�~��1 J��n�4�L/��\�Ge��8�i��8u�Ź��ײ�}�v�u�`�{6QZ�a �����N��Ѹ͊��U��(�H��=�b>���-y0Oƌ��'�xZf2yfzx����R<ݶ<<(�����e�X5ҫ/�$A� H�����˲�N,���qك��\�H�Q�8��ߩ�?���Pu�w"�ɘ�XIU�'�u��l���	ּCĩ���>���o@�"����F:^cyV�8�\�U�YM��>OB��q�Y���SQ"G�c��)�PvΥ�C����:������y!ʁ�ʳ4Z#�3~to֪�6V�x%�s���숑6�ol���syK�k�!T.��Ý�*�.��t�)��~
^���2a�n��*O Y��&�B�[�[ٙ�z�_Ј:��~�ߜu�,��Y���&R|���7�Bg�����}���M��g�K=_A�HX�uQR6ۏ�x}�����x��!hj/��h=��H�^�'��=S\�t�KIK��*)����D����E�V��X��� #1 /���{p����-n�~e��b.��2�Ef1t�*�����'�EG�L��E���[
��<�߶�ZV:�m!�
|bmf�<u
>���"�m\QI�by(?H9CT���2�`i��J(�)F��ȸ�!�8�k���v���mB���_F`���W`���u��{**�\�0��t�ٟ�T��	otZe9Y���蚈qg�����G�ct��Mީ��WOh���[�B��vm�N��iʜ������C�zw��}ۀ�ߴ3����Z5[Q�ڑ�wϐ�t�M�[��3.u1��m�!F�yr+)<�'D��̦ѯ͇Jx�+1�i�(�p��~�G��:�I��O�� D��%X��*�{;g���VL��B�^޸�k��yԔ�&�s�����G$�1�HN(ӎe�ӌ��gĥ~4�Z{<藦Nr��`(RGf��|%�yHU�� ~��UY���HҎ��k�hUb�oF[���T�ɗ2��C&W[�D�t\�?�����"?CpEp=����`A.��n?sQ����@�`�E�6#n��+ܓ�k4���4n��-1�}�r���FEg�Ӗ�1��e��f�,�kG3�ƶ�PL�u���b�jT�!K���6�a��*`�!m�%|K��u5�P*�T�ڲx���r��C_���
Y�Wʷ�W���7�e���dŻ�sr�l�(ye�n���ҥz�JJ��v�~(��H����t1h��-��xܲ�����#���v�y�H�GCO�T�tw����%\�0��)��q�sn�ௐC����g���Pѭ/a$� _Nx`Jͯ5i8��_u�H8�	Ryy�=��|��0�Ŵ��v˯R�M�\�J�`�N����u���A �wi�#ã���6h�z��y��ZJ��@�	�M��H�|��X� R���ﹾ`d���H�^�4*f����"�j��I8�1
��O�0�?o���8�b������ʏ~.�Q �&5"�0�Z8G�O��K�����v�sQr�{�b���ʣ��NPCD�n�;8���gI)������i�Ǚ��L=3��#�{�$��TWY��b^��r��
�lA��aza�ZS���`�S�������������b%z<U~����Kh�B�t��\��HV��m�
��p2kwl�s/b�~�Vqi3��d���:��E�6�z����Hw�)x__�B�\�V8�|�	n�ٳ�Po����ZA܂���b��#�q�<���hq��%E���H³w�����=��(�ϡ���N���ի�]5����y8�JW>��y���QW����D�fwNeZA���x�F}�u%�EL����5X]]KHU�8������(�80)�Z�Y�;l��������Ö�
�����GoE�ʳv����-�%�漚������Y
'�C��ے��p~�ִ�ϕ2������	����C�V�ŝY��>��b{��C12�㠔#N�7�m/��k6<� (�ڙ.8�s���������}t��Y؟��A��1�R�.j��I�q�̳��J3���j��D�""��ڂ=��	ζ:�gg~���e5������l���At'�z�z�X.�����/��D@"��hY�G>�k3�OVQ˫� �o���z��@y�6΂	(���D�����RC��j�q?i�$�Ua�M���_�?!#�ވN��ʟ��#���O*Ū�U�B*�a4)D����+��1�jf�=�M���躶����Q��]GW�	�%�*�{��ܝ�u�ٰF׸�t�
�v!'?}�ޘ��kZߧ�
L��\KN
6�`gB���a�y���!d�� F@+B�mv��2��o�f�Ք�ڸe�0�2���֐kJ�6%.'�	g��C�Vw���	,4s��G[ߴ�4HC�%���-�������6�e\`jX-*0=B4R#�AĔ��Z����J�X��٣��Ͽ&We�+a�9m��4�t3�ߺ��\�)b���������]B+o~ܘ�@,��:�Ř��u��@�*��o*[HP"H�)&�=��o������:
�_q�� �expӛso�g�އg��	/`v�n^o;	���?��sj�Q�1��� ��w�b��+�����yNE��WR�o�v��Ou�^ �1�H����_�A6�r3T�&�$5rQ�OYS5�fY��̧�y.D��*�ʮ�d|l=q�P�9l�|&��*6�d0C���:��]O��0�sBt�cI^�`n�@&\��iL ��`qY��r�e�%�R�l��a��"؝-G�͚�#n�府pd@8f���jky��ˎ�l���E�Жi#�ʂ�rr�׿��U�7s�
����Y��9���l7[@��42�F��~�����m�`�,������@y�h5�t@�ʥQw�>.c��E���!
�1��V&R�j(ǩ�w?�^|��nK�n�hlF�����W�����Hr�\H�y9ʈc�X�����\���j������}3u���m!�d�;����?��sq���{�H������p��������[�+Ɇ�NR���x�g1/e�7(��0�	/F�,j���E�r4�ݦ�#��I}�5�NΑGҩ�._���w�}�`�ke&!�+����� ��gvo���0���Nw�����Ӿ`a��җ��9VpA9[!�ˁ�@�9;����Q��-�P`�ވT*�5��Z���0�h-r5N��� �jǴ���篭S`0�m��3,�!���/��}0�^����͜q�I��U�q��d{���E��c'�W��D�yac��[\�D�� �0w�\zɈ6�µ����Lbo�,�s�f�)�%{TpWV�1d�=K�^ƒ0aD��&��/5/������7&��b�Sϟ���9�t*�l�B\O����k��S�݋s\(���>#<(���v&5\���/��-r��p���(dY�J�V����]*&T2�5X��v��Ĩ���dR�al��B�S�U�׋�KIca�!����K?'�W���_�����_I�BA��1�������w.�ܘ������B� d�J��L��P<��t��o�2�bZ�]�ELHj]ZԠ�ޭ�z�c��(���=��\^0��k ̅������*�F#c?L����ב�I�]#}.]�j��t�4�j��65��0TfQ"+��0I4l�x��o�X*V6�և.��f)͸c$C@_��,s��ng����M��{�nM�{I�K�*�w�R��)$���d�Sw�K_�?Ǔ�O�6�(0B�|�����`�� ~U��d��D�;�'�Ș�
h�~����}�v�6Rd����]�	�0���>E��ּS���Y��H�pTU��3Eθ�����F��I�"�b���5S�ʊ7���!��ΤHa�A�ޮ��:����H���"��Z���aG��D�1�cR�C<��9����g�6EB�C�E�1Әe��X�甸�_�����b�9��ٰ<Df���!a�f���@���󀢅����7���~j�}\�ֻi�QQ^[!�~>��9���tm�F��/�Q���Fr-w�k���J�+��4���P�Q2�8F�lY��GF7�._�����'�Y���>�������F3�X����?8�&�A�u��[_���v�RFUjb�㾻��<a�3�S,�|j��b�����6�h?��&Z;X�k0���
`�wЙ�Q�rɞM�4*h�[Z������G�z�N�%[����r��3����/Ԏ�`J��K>C�/}DX�+���"�c�)��Z���V��s��EL�z�9�ys�顿b	`�[fTz��)�cm,J#Y�{�}!��-�1^��K���Z'^K��`����F��'��̝IZrP-/F�C���bʱE(�a\M��8��Z94�fe�J���t��_�#X��_R���s�����W�[�!���-�[�7U����7�j��X�9c�e|�q<���W�Ѣ�	��":̟y�*@O4�,AD��5I3W���. #�5���IP�{L�R�*�j����2M�S�YbIB�Nn1%բMů��ťz��7�0N�Hi�D�P�_�,J�{� ��3�v�y ̧^P��c��$S�vB����aB��'�E�r[�w�Jr��:�h��Ő�����x��tPZ�	�.�G���`�v�p^�W�ʃ��F4��!&m��^2}�{?��^��Z��t�kx�YU�/�l�^9�*��]�?q{����imEE��G��YHKd����&���ߗ�wx��S,���s�>�}��.�أ�H�l���N���{=�|� D��<���?�K���1\�9�TUK� �����H�e*��%n��)�8��k�,d��� �A�X�Z�y�w���~�����+&� ���K�Cm� �@�'���d��v���I���'�*07v�*l��$�71�Ϡ$
��qԌ���cI���k`5ğ6�AId���F�H����¯��IԓC0��W����p:�����Q�l{�:��)�� �k�^c@�������W��{|��9JrG6��n;iu��`/=��f8�a�G&~ЉR��/w�������,2�T��z�c��cq�9��1�-������(ĒI$*h
��qp���O�P�ڕN�"TJ~)�`nb>�	�_`j��54N�hpo���韕޴�N�$�a��ƭI~7su��\5�b�eE9�8��)����Hۿ:�Zҥ!s��ŏ������L���Ӏ�)��Ѯ����+|��F�LE� �vB%�k~��:�2�:[G��3��w�%7������k�~/��3�{5�G����S�-Ur���<��yKd���ɻ!��sދP��_�Ч�Q�o��G���<�'�e�S$�"Kʖ��s�=k���<��W�%G�ڟa���l�ϦD
��5��ؒ C�{�W��
22'u�\�9��prGd�&����^]����k�D�u'���F���=2N:;<ْܻl�D�%�Ww7�2��L9\ט�V3���;�O�Gr���F�
��;��I����A��:{���j�h�O��0mlr2�A�{3f"�חR����=���8���bHy@C <`lM��!%ß������-��� �;����;���"b{8��u
;婅L�P0��(՟��<���,fC#�Gg"`��=�)������;qU�GD�0�"���f�0�B�´�,p�YǸ��^��<�9v�2[.4�13@�HX���˨�Ҟ��D�9���O����"�:K�W0[r&���.?{h��k�I��ӴT���,&�����(��	Au�bڶ�v�l?�`mz��do�W��ȍ����Nq\��U�A��RlWP�d�8�נ�u 7R;j���d[X�����Of�6f`�s��Wa1�1k	9=�~?=h��W�;�3�W���*��!(�%�O%ݒύ�#��,'��ߕ'pxξj�9  [<8�/��o�NL����J e��PcM�g_
��`N"����_�~UJY5�68���]���2�.S#Y���z�ce�0��d��JBPX�����D�E���q5�c���Us�]�i|�|{�׫*�p�݋!�5��;q~�� �,���\�&D�7�.�M�8{�)��7��SJ�`��&Q��|k��Mj5x�[kne�Ʃ*E��&��"u?�䑎%�N������'�m%�$Uh-P���{6[�8k^��O_{�9���V�b���K�f����������c+Vl�v���4���10F����N�	'w��}�0������GD%�ie�]��ӧ*�
�o97o%�|�����J(W������"�5 �h��鶂MU1K�ͤ�I;F*�{+��(b�∡�A�kpV�ty�4-� =ʗ�k�����N����N�|#.h�i�-oh�؃��*M�V-6Աk�ֹq�P�9�<v�-E�6Z���YIV��0�&�4zU�����_]�y1�� ��8��g����伊z�s*���[�Ci�+�n/��v������R��ɿ�����+�{GA��=�0ԊK��>@�^��2C��E�z&6.P��J��!���a�l�tƈ�լ�F��:	��(Щ�ɼcd�<�;��i ?t��QdW�f��"8�y�"��Ȼ���8`I�I��;���c��N��1��e�h���ʺ�H��}b6���b�����e�f�A�LR�ֹ_��%�Z[XC���~�G���ҝ��Y�C���Ӡ	����/�M/�M�Z���1�=�˓KP��ۖ4�)bw��_�����\��`~넃��u�+���$	��\Z˼I��Rz�-�ŝVXdؕm����l��_V���S�;���m��#����΢~{�.rѕ�0�G
�9כ�`�E���Hp�4ɛP�S{�.ٳ�˵���rb������	vZ�ѩ��Ѣ)P�c;�l�����F�+|�4�R���"�Փ��K7/iOR����3�%Z��9�8��5������/Vz(�U�S�aX�<+ݵ��cW�E��l�4X�����?�s�Σ�u�n}��	��g1A]i�����[S$�>�`K�II}����?"��׬@�.�X�[��V��*p�K<i�!B�����V��/�F��lA�-� �֙q(L�E�V��,��*���:5�l�?]�г�s�>�l�׀_=:u�4_���h�[��,��Y�2�+Bi
C�-��0�OWU�,���!(��>v����k\s�<4g�ӆ�+�)�*`�-�a�t��T�@�Y�c�IB�!n(����y
|Y�P����c�5?V���g�Cg\Pl+.^�j�"�I;�-�D��?D/��tP�8"H�pg��u=~�k�%˩�I�ݾ����]����~����&���@C���D.��[����$U"J�J1����ЂB$@����ê:���R5J�L]�AH���d�X�\�S:�1X�qlv��"�(>�CB ��A�RuC�{�i�njPW(������ٸi������c��N�0p�L��~�)�/
��""ԋ�.WK7�r�D�%���g��q���G8)듕��ܥ��f�p���?^Sb���r;9��g�.�yZ�3>�kL�}/�B��_B���q�4)�$	��a���2qI�A֖�h���Sg壻K¼6r�E���]X"��U:+G߸����3yΈ���U�(��u�K��� *��=�!%�S,`庀�j�6}������c��.������Bcl"�ϖ�v�|�Qu�#�{�7|C�-b���q�M�����R`i���P��$�@���c6�͙T��4g15#&��ʖ.`����%��	����/��+s
�����.@��}&�7�#��a:�(���ڰ1H���֨#Ɣ�0��i3���-���_�ps���h�x��PU@FH"����мM_bP�Ʃp�ٕo ��$�4_��čX�E�~]�W�{�������3����c�(�3j?�����1X5�?6�>�ּ'[��o�q�YT�9w��4�)����������6o�˺#v 9Ѳ�\o�����W�"��^�Ӿ��ck����S�
Sϙh5�8x��ed5ɕ�\#�V���J+�ջ�cԮ�a"�[Fy�7Z�ls��mbkoET�g>gqN�0J�m��1��@��Fv���I�� �j֡�A���o�t{% ���~s̭�s�l")���׳��9R⸥�D�y<6���w��;�S����T���}�p؎�ϐ���(�kdn�V+_��nl�3�b�ll�6$��V�K7�`N���E��2M��w���xxa?Dڡyr«�?��f�|��i�!�wT�t�7���_|�g_m@q����]+������;b�I.
]y2<�e'o.����Hf���}F0��^�WR^�,�"����_�EP<�S��wK?�����z�~/���:�]g%�^IC�x�����e�e��]��������1�l��2�k������w�v��ˁ~�8y{�O�Z�B%����N�QW�������Y����/�#{=��&=5�o,����pu���m��V*<��mں�<?� ���0(�8 }������]�Ѽ�5
?�x�/q��9VYD��ĐY5L�����X�������|��{LM窣^�R�Ӈ�|f�~��#�?�κ�^�>������e�z���-T��� �5ᰯ���v��&L>�-(8��;�s2S�l(��t ����Ta��ٰZ��P��Md7�G�bJ�+�B��NV��]�^�3d~�cYߤ�z�2F]k�.���ג�����v�}��r��0�ɮ=fP�^nk�)�L#�e�[��/����[eV��z���7��4o*�:o�οk��1��1�}i>8��h�C�� �Dԅ�o皆���#�$l�'���OP9��	��@�f�����i� �-`��B�c�(���� �8J�%���G�Od�Z�/��Eʚ;f]�݀�(UD�	mz�q����C��si�n3X56_3��>��o�A����B|~/�Q��r����Q�.�0�f��֛��v�f��r^C%�%R/6}�k;���+���<yYn��0��Hb�䟰���TG#;2uP���݈}y��zAT�+�s	�xT���㈨U���L�_&~�-x�z4N�v�����߂f#Bݲ���"��[��p�?�s�a+�gJ.�J�aϛ�<����V�'K6����i+����R�o6�ITr`ނ�qϵ�YS������ۙ��~���ν����Q�;T�'�9�����K!Z��O��D�q-�%��q^�/.�V� !Cۺ噸����?y���r�`G�� ���L	��]e���77#�,;9)<1�ғ�X��Q���a�뻿���:�$�� �Qm�sS,]��":��B�7g��Y�;C���{8z@�[�	�}�3�؟0��A�E#4�	]J}�`w�w8��Y[�{��[��۾��}�2����X�<�*�&�<!�!o���N��"�[pYҠ]���hc��>g�0� ��M}G��c4.3�h$���ʌ^���)��Иm����46D��Ο�d����)&9�(%������>�UJ���Uj�0J<�_N�����n��9�bCE�N�fj��B�˭�	��W��ʀ�XCH�BU�J���j�N����p���*�j���'Z�#t�,�^��W���V#�>ڼLF�	(}�)}G��=�M�s��9����V����e"É���gx�B�k0��Ū��4�|�}`�5 ]Qڂ�W�P���3P�X�@A���>!��Ef���|���/��������l��\�&���T�?c���%�Dha\��y,W�"&��	F ,�b���3F�Q!����nZ\[D� ݰ�^Wdb�L��Y�v��Zh}�ϱ"� ��o��ɥ&�3lV�����W��D�d�a��-�Oq}Ś�G��(<1�,2�u��Bذn���8��e����nj(�T;?�����ύhBd`h_e��<��Z�YD���� f�D�Dx~PnX<j����"��<�F`d����f�����r��l��?6v���j4{��B!�'~j6��UÆ3m�,b`���U,#�"�7BP�{���`����um��X��N�/�F�{�KX{r�\��"�K�{������My�UG�|��ӴN��Ԩ�m��3�W��#��2#FDLB۬D���ݝ:�܇P���6�UO�K��}v��{g�q�-Ur$�&Pv���+�K��j��[�I{�с��ֻ�8+�r��e,R7H��3��g�{�'LK�
�Z�$392��*X+���o޾�(�6�������'���]�P`��(LY�"���N)!��ޢ�"G������(BrZ���۩�\���cb�韵����q�9�Z�x�`�`nw�����V`	A����g#�� �)f���m �2�����c++���i��E�O�x�o1T�>;�XX�����R�3�Z�G�=�{�)JMD:џQ�˽�S ��ц5���9�L!�l��-�hP��5V��
�w ��ͣ@AdZ;��P�(��eD�h��I��S�,-��wh��Pg;�2�YĎ���{�������P��͌������'�#�|�eO[��՘�����]8��ѯ�zs���+�<x	�he4bU�RUM�19���<��at���S�?6	�<9h���=>4��g2zPC,=��xz���h���E��U��Hb���c����Dv�����̽��?��bH4С�v��l�!)��h��+��J˃�*�]���;&����a���^%M˳�h��\9}�e3� 7�U%�ϫ�Iu�8��'OZ{�* �&��o���f����g	� �_�@��w�%�~d��E/P� �K��X��4��r���[bIi'��Y���Ο�~ O�̋�!�~xd�
!Y:��"�׵B�%�vڰz����tS7/�����E9�m�����y���"��o���G��0(�2�L��LЕ22襡E�*�-���m�öS�Ve8$�p
%���R ��~y҂-��FT������R�vQ�19).�<Wގ��W��?�iA����!�x�jSeS�lO>X���v 挮̘5�Z�2yK�a9��ԓ@$�ڢR�i��k�vh���5>�`�LkOL�3#�	'��g`��:�˔%:��~!��&Cm`u��6�08[���z�[���}sz��~��g���qS�[(��5���'8�W�&�q�}k�s�p��C�/7H}A�fmD��I�-6���ar�tfʻ�DKٍ��_��3�V�e �1ܼ��a��Ar�X,:
ރ��%�[��ؑ��^� Bl�P������	;�h�e�e'��T�g�+��lx���TP����@�t�����Ms�-�Ĕ�S�������*vJx��p��-Zķ�u�L��z�n����&�q95�F7 U�DZ��
��"�C�Q1	�w��1�@Ѭ'�{"�
�i���)����x3��m3H[պ��4�K��$����=���ĺ�`��kǪ�3����f�<T�lD��]	��g�����A�S�rB�{}kP�f�"&�O����7��;����_X4B�x�\-0p�-@
�n����y4 �7p��6��g��X?�C��������F��:É����oX�
!�ќ+�b�8���j�(I]e���⃎H`ƸfM��S�g˯)N�l*�o~M��� s�U��	R5���a��E�b�c�)�U��>�T�>��D��g?�֔�v���P5P�"��Z�Z�W��v:q�k�2p���zA�ƍ�>9��-�IC�Ϩ�i�2��P���d�n�1cNi������o%�I4���=D'l)"6�R���Ĉw�~{����>5&M�GP)����Q0h�c��?��I�ŧ�)���r{d�U�;rS�q���Վ��o��
�?h�� ��z*5�E�'�U��R���%P-9=���M�x���m�R�e����~7%$f��rQ"&jq���N�X}�� PT��dz!�@Oq��r3�7u�lOG?��rL�H�c�a��Bl�:���S� L�)��*��h9e�J��M�Tj��@���p[У�E	,����]Ֆ��n�Wr	�?�z�A�~ !m��{���\��a�O�u:�hXK��#�z�Yk}f儦��8������d�Eq��`U�{�,!c�n�c�ɑϵ��J�K�	�Χ�u����n:��K���dw!'6���� ���%?��9j�"a�3s��"0�St�$L>�����^�Nv�F�uX�Bm��Κѩ�V������7�����٠q?�yF
�D"2��,|߂$l�w�|Y�����U-�����Ј��*��h6�������	�'���Q0���P���uЬ��d�p�+�~��U%�+����������m��<�Ӄ������f�&�d6=�� �S=�B]�߲�����'Q ��P�n��߫�`�V�T��嫴��{�[-$�٫7�".�!p;���QY�Ur�Pe�Z��J�������\�5#��s{�Wy�Dk��y�Sg@��v����a2��B �T��4l��Y�~��L��d?�A�~���[��{��'�S��E�����t7��5�^��ƍ%��s ��ی��p1�2[�O1m�i��-`<-��PD�G=Jp"RY��T�:�~3��a�V�
u*?I����w�i�������BQ���&-$x���m
�ħ��[5ZX��F�ƤKa=�1Y��Kp�)���[����W�I ؤ�b(���0EX��eV�΂��&�5���ƪ!�������}u����{(Lȩ��K��k�`�ߴ����1.��.W�4y�F�p�M�F���0�c�I)�n����u��a�+�"�� -�Ɖ�Wa���#t�%���ˑ|0�VX��s�|��d�
� '
;$8�W:��P�J8���Mq5�~���]ބ����/�S��.����>��:�g�shߕ�<�k�ݚ������b����}'*�s���������s4����
c3TkQhAS5�P�5!M��?^�k�J��Лg�p��2���@8���硔����=N#,F�l�o,Oz���;Y�jX��\�cj�QϘ���Q�g�\�L(�26o�x�J͸�����ie��ɮ|�9~��:	�J�!H����8b`O��I=D/j� ֛�o�:�c�<��\�<�(_ �c���=� �N�����2��&wig�m�p��Fכ�b :8��PzX�P�-���Z��X�a��o:���2#�i>>�,��UZ`�	3��:�/k9r{4S�r���Uݱr3��L��\L���S<����hV���3�=䯚�71��Dz�}�oE����˃����-��|�6{�������Y�t̒O����W^�^M�X��R����m+��&h��R>2[U�&��1G�Y V����U7ل.^A;ĳ���*�MʲP�#z�I�H^E����&M���F�E̥'��pto�
�~���l��|��R�g]���!��\T�T�M-���x�Y���h���D�r#짶��{�ծ�'&�_>`5����f�0��;�.
����`��e��V)� �vVrM(Sq�JW����y�?*͆��8��l�J�ٝÁ����1�H��P\�L��x@J��ܱ5	i(5�Ӯ~7�22q٭����rUA��a�d'HHY���kZh�P��ݶ	s��b ���-�YĊ��>�/|J�@؊�J�D�!g�%S���2K�M�uݒ����.���o�h���Lד��Mx�z����Q�Ђ�7&���ޖ�0Kp,�մ��Qv4�h8�=��b�H�k��.�nf�0��׳�vĪk&���L?�J�A2F{�[���T9r��4	}��#W{�"B�~K%/�{nq��¶���� ���V ���D�=�$d�����l}v@d��:��t���1d
���SK&�	wO�el�-���g����ǚ[�i���-ڦ]�@:Х�L�7c"0��#k���j�LUX�'?�����I}\�h`������w��Y��/n�`��KÄa�>�5��F1���N��]@���qw)���mi`�o�_,��I�F_L[4n�.ޔ���'��:��Z;�xw��uTW^�����t=�${�D������Y���'�T}! �I+�<��C�\7���HE�Ӷ��"IRS�l(�@A��p�n�o�� ٝ��A��M�5^�%��lKn����p���s���yKj��8���2 ��!_��_��� f.9��v�O7���ڤ���D�.%��t�U�����a����mg�����ҮcS� ����]�Ԫ�4onừo�9my��7��_/��uPߝ���������KJ��M��B4���>�I�?�ͯ�0��jBY^���7i�" �&��|ۼf�`��g��X�{
���+k��MM&C�@���M6ntBʔFѹ+�Dh�L��ᾼ��#��B�*��m�G��߼�����4��i �-��M!.�VVY�,�JĢ�o�Z�y6���wz�+y�u}�jo	�F�B�sDq���ÄF��Y��q�"��tP�p���ϋ��uze�(��<1(r �ښ3���3�,�ҶE�A�����zVb��s5=_|.��s�)��ןg�m2v����G,6^i�yb:+�3h^�Çq�8˜�#�߻����O����� J�$�Җ�^PT��6vɟ�u~K�v&��bSѴJW�Z�~klW;r�=yq?X�ԙ�+2jf&�kĺ����Z*Iy�b!W��o!����
*�&ht2e�,�?���X�㈩�m@�����jr�6L�\����d�9��{�hN;�Ü�����,�%�6�1fB��+�2�l��g�α�����J� Y���m�<�I߫B���\݇�z�+?��6����a�D��b7Fkރ��M�gX�u����ȵ�hP<��}�fLh2Ά��ϯ��JE�Z�F�9Z�,xpҟ��c��g86���I&�ZPm�.!�i�X熩���k�6�w�>�&Qx���ʾ�4�7�(U�VjA��>�p���߈�pO�)U��nh�/#$}�V8eDL㇒"��r�� �&㥶фis�͓��T;���<�VUp+C`,O��u[����Mb&'0��\��FO��g��
������r�4�ԚpK�B��Lu�c�ƚMwl�V��G�s�B�|�WI`P���K�R�_�^]=J��!پFHs<�'�m�F\�x'D��#�����E.?�g�'p�\� �Mu�2f[^ő�����.�A=[u^�`�)��&kj�H�D��y��&L�ۆ����ĖkE=Y-v�)�ƥ5�ĳ"��3���I9,�%'h�Qj_� �Zz/�@��k�Xd��)0�k2�x��C�i�=���lf�1L�T#�.4Q>;=	o5`lc��n�kL�,̧ة�ʦ��߻=�����H����p/[yd�&sH��{�I4�����DrcU��$�����g�_�QP ���X��s+hBv;X�:��t �/R��η��^�dυ�OL3����e�Pu\2�J�SD��j�(���o���+���O��z��xG�̘R(�A�`�{1�i�bzd���1��
SX&�}�P�W� �V5�٢��^7M�kLK���#�|�і�A�5�jه3��rZ�a��@r b�����V@��QV�M�:��)u�Z�ڮ��S��}H��ae E�k\�v�M�(��zZ��mxe�<!�e�V�A�Ezk�Q�)-�o2��h-+����_17���:0�_���/6��b�j���BfA+]��z1T��Y���IQ�O�2�~��8_&U_����b���z EH'۹�>���g��& Ps 3|B���Ր��������+�vm�EPn�W]/�"̶i�[N�����BVW%mO���0����2#T9���]uU���rOϴ	�1�ŧ�c3�����{�s�j�wm���r2}�鬔���*^��-�+w��侪�����ٙ��:��Yta5fHȾx�����Q'�B8�>�)Mh���ϓk�DT��spwP��x�3�a ����h���J����͹��{��Ϛ�'煜�"xM��Ak�Zά������ ��^� "5gVFė�fꠂ�	����v��� ���C={�T!��X5�+����Cވ&�xN�Y3�l����"'��L)���JW����l�9��U8���[9+� gc���f*��c|�o+�٠xYԱ8,�}���g����h�#�!��Ѿ.=��%t��ɪ@�?����-ðULc�Ë��@8��4:��t�jv����9�]0Z��W�'�Ɔ
|S)��Cʷ�{͋�临/�l�ri>�A��R;�6�i�[D�5*���%[�ma�U��	��~�}��"I��6�w,Z��]�>۔5sR�|��nl��T���̢����s�ߜEq�*���@��z><z.����*32��'i��U�b�! �	�P:���ͯ~�c�d_�-D��� =������F-ikCë�hψ��q�R'�ƃ�#�"�N?|X+��P�T7c�O����;,/<���Ā�+u��e�I������>���Y*
/BX�AȄ�㒛2d��pgG�R�>a<M�H�\�;<����V����WjغJ,i�`{�?�zE[���8���~䌁�|h��pt�(j�W�1�����Sp���*��c�d	�7�ưy�%F�5���-�_�x���Ě�}�RE4ľ}m�R��x���� ���4�'u$�wu'}`�p�SQ��H�b1��� C�L��A`b�A|��=7x��`ԣ! r�8� ��Q�D�8���T�u~/��l{�>o�O�	����"W����Xxݥ��+���F�{IGџ����,g�zڴ�`c=\A��fu��?�~=�^�r���ݭ5�Q��"��~wz`�J�� �>7%�>�^�yd�<W��KؐP[��Y�%җ[�ɗ��m��Ɓ�1P9�0������o+�ɣ�00��
��E3T����QF�~������3�voIp�ꂓ8w;E|p1�D��jϘ��Nz�Z8�>1�9y�K��Lh�3��a���gM �@[�.pc�����LF/�3�,����0̨�TYC��$�+�We��}twZH"�P�\�`�UКNᢤI�Ln�sdW��Y�'b*�S��{i����^M�P����:7�ax�R��2�و��iT�~cc$K!����ܿB��Wo5�5�>í]����^��;��L��q������� f{�1LA��1B��T��޲��A�������E򐹰��+���Co�P�j�v0�ŷx�\�fyQ����_�l����kg*�ct��p	�㏋��Xc��������1åal�Bh��G�m�`I��3�=�q�Rz�+%��HJ�&+�Vb~�]��>��DT��?CK��w��Y%�~�s~	�pLڎ��Qٲ'6�����6#������a�Ÿ�܋͈��l�x���<��Nj�/�^�����\��N4I]�{9q�t%,cw/�_�	&���5��<�v��1	!�E2NO=L�����L=RZ�-�����I[9G�ʮhm�m����$q�Ң� ���3bع��1�僃�9���\p&��&��}��}U�֣�dEt8;�/��Gi��*�zL��5?��:v�"�_pJ��2��J��I�0}@�*L���3m��;[����Q�M�ķ�1ҹ�k�ݛ�B9��ƨ�N#�ڜ�3T�z�-㨆!Y��N5d�O?!�s��}hh�Y{��TBH�e����ksA��"���m�����\?I��ߛ3QUE"T��ٸt��BZg37w��E�J��p�'����^��A�s�s;�W:�Þ?n�T鰫��ڠ(�����nI�&�'�ͷ�g([��CP���Y�^���t�nõ�}��8�H��� �x����Jܕt_..�<e+�jխ,��}�*�a5�@���R>����ٙ�����b�%t��VGqI�d��xg!=���x����F���W�:�,И�RN)E��rUq������Q-�F[A���ѽ>�r�vu�t���?� ����J������J	E�$�9��\�4�t�T	�߃� g[>��<==/6���_����_chu,S�rIݲ�ֈOԍS�����4���
 P
ƃ�h~,�58%�@:A�"��5M�/��:宱p{��`�R�ӝI�y[ҥ�D�3#���;�Q���F����X�r5
�#��e�_2�Y�*�Q@�2�����rx@D�j���I.���h������R��C6��	;[@2�d�RH��'��S�z�6���Q7����b� ɵB�U��0W��A�S4�������$��H#�(�((��L�4+E��LF}.$���>|F~A�u(�#��E)�O�l�.g4��Si��3��>>�T���1Q�L�9ѡ�b�����tG����r'�γ-1s��Ͽ�V멧62��Q��WS�|ER;#-�G��F��_�ɫ��-��r�.c�E� �.�w�-��(1��W��;�hV<���pp�T%�G��iޕm�OR��
��פ0o�A"��(E;� ��t���� �|j�9_}�o��CT7�.��h���֘W�]��[��g�C���{ӝ�&f� x�V��_����j�����dW�u8@ζ�kf���Z_Y�g��c�@�%>�6���n����˴��$��C�M���tuJf=��؟
��uh��2C�GwH�BP���L�HE�뢯��Q��Q&6�ep�^����Xc��
.sV�bV�C/�~B���Hv�K�����p6���:�bf�d�X�
ߪK��GP&�7����u e��!������v����:�E��W�n����ͷUd��
pC2�&�+�o#�h�n�{Đ�kf��tCI��Y��6��/�$h+�Rb���?挜�y,v@�e������s�w���������CR -ݔ}�W��`JJ�5��������l��g5�4�C@ ���ϓ�j