��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4B�#q�@�;<t��:�[-���&��5/(���{���i�9�о=�%}�~BW.p~+`�l�`��c�����eB0���iأ��䧽�|��b�E��bK�����P�Chw��ަ(�!)������OH��}:�����>b%�7�dH�^��UdS1RLS������i��k0������[����_�:���b��Pv��&n�t�23�1�i��LF��m%&�X�;�A��#�M�L�#�b��O���9c���q��4�1�����$�4�/���mס��TT1�ߊ��7���*��AG����f���s���lc˛�F�/�qE�����5]⌛���F�I�7r�rh���Jd�����:������fDȊ}��{�����p�k���/c�>x�׳ɃG|�PQ��~�R��``�������絨�9��x��:$�I����S�p�_$>*_�W3�#d��f���rB���GR��m$�'O�}�qbY�e�iWk��$�>4paB^�,�������?�>�_r��i�Mע�6��ө����U�`�Y����$Mo������%w������'�٩t�c.%�����`��>_��� F��"X�>H�g�C�D�����v�áA�m<C15ЂW;A���Tk[����آ��ݻ�ӂp�����b� �Z��E�.4B�Ui�x+"����;p
��(�e�G�3K��02�����&zl%�;RXkF:+�ŒҞ���7��'ã�+6_��5AV'c��ߨ�/͚��~e��wc���ݡ!�l���}J�[��P�����fC�］km^��I9���Y��r&�?dUy�����:��ݻL��p(��br��L�f�w�$ر�5j��M�>������r���8�(`�*�Y �@���'ӗ�Y�"d�lU�@mu��=���$~� �\{gm�ٙP��� ��������wx�(\nQ�Q�� ˯o �Zv-�o�ʬ]�&�7T�X:�~ʣs�G_�rF":�o"Y�0�g���1��,���j�(R�ڦ"2l ��������t�QΌԀ`/c��U�Y��{q�Ұ���.1�ün[���0d��jL؃�
F�'��!�3���CnN��0�V����5��<|`%K$H3=��OPb�#z�>��S1�^"IjUD���+���R��o�U6��4%%������&]_݈�C��a�\��7�3��C#!��ՊX�D7ܓ0�yT�Q������(Ώ<�_3�ڰSy��.X������N�ն�1�.�^�	no_�J��g��/�s"�LY�L��>q�$r�q��9l�ō��w��y�|�6+��J�τG����'��/�
���Y�ڸ��?����������¤���P�	���8�4c8�Z�~�9��dզwJ��35���`s��		�eb&�(p�@R?��I�x.f�}No�΄!�R5M��8�l�p��]$��]��?�d`��#\�X,�4��ũ�[vme�S�B�X�Sj6���9�&'D�z�O��Ŷ�B�e2W6W��Eo�Dby����4�� ���r;����?�@	�1U:�P4q]�����p��x5�rm���9Ԍa/-BV�'�!B:�:@ ��Sݍo?�ƺ&[D��=�5N�r �R�@������퍅���/���h?��٪H����v�luE䊐e����T���͔�L�Z7O洒:��E�I�H�U�E"fp��+_� X�2����/��-98jL��VɎk�:�>ű^P����p�x�
�(��,�%8L�g��
��h��R���"��sֺ�����zx�y��rQT�҈�R,��Z��Y��2 ��������3�N�Μ�������yxv�ꖝi�iQ��5��8R\ X[�@u�ws�����85p �r$��`�O{�q���-���b`9'#0^�RG�:/ d�ы�m1zi���@���#G�>�&@]�1r�eIRb�u��)��c��p�+)wm��{��Iy�O��GO^�6�B�`&Bw˥����ɐymc"�Kg�i3~�a`��:�G?s���4![,�16T�@�S0_��Bz^S���8�<f�p��'��%����:*`d�@G&�Уn�/�C�����<on�a��������x�
P��ْ8�J���扅K�ķ�� w����~6`���w��"$AHm�'6M�5�a<�[�I�T�������}�E�� 0��C�f\�[$���KM����?b�#+��z� >�:����[p[7��8!�r����f���ڭЈb[����ϧ��������vx�5M��f�"����1�vsc3+Ru�7�]����7"��+�[ >v+)�df�!����D�.����a5�dj�5���s�2
miK��<V2G.�
���]uf��z�Se��"��1%�!!��n�E��{��2Z)'��{rE�xK��Oئ��|�*1rj�6��o���sj7;�&ŵ�ݡW��Ot)A�6}������C'8<@	 ��7##T��U�]!�U�Z6��j��[��j�hߨcH[��KovY��>�Y��+������2lGtka�a(X����v
,E�����Rq���a�U��%Rs���������Ҁ�4M���F��W����[�`\��@Dh��k�,׬����+#M��1ķlRܼ�5>�H�:r��]*n�]Ow)
��W6$w;f�~��S���K~��x۽u�ؕ��_'2O?(�3���z�6�a�޵S�f�e}�
�\+�||�W�H|�:Ih�.�<���S�����7�ʒoٽ�<�DG%��n���`�]�n�$����h�6�Ҳ�`��\���P�̿��A��?�JFL2P��+Q�oca({/l��b�o�*C���X$���̎�X�v�ظp���i<1�vf5��ݯqN���R0{>��p�Xq-x�`L�5s��)|P�Ԟ��0,w�"'/
���n��r������Ho��N��bI�3�