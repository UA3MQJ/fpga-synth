��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su(�}&c�A������-A�*{���G���ٖ�� ���OЖ��rf�Z ����j����̑`�֐��()��=��Plt4�p2r������Z �J��H`��@p��k�f"<�s
͔4�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��։�������7��x�y]��ѬIf-fd	x�|���!FR�?XG�G ��s�����R)����Ƶ�G���Ex��E�f5�`E�m�4���Ƈ[��dЃ�M�`h��@}[�k`��W�&��RRI3� 7�Pu���~�X_�Fh'��m�]to���p��'��ż@�
P�%���"T�'Hg�'���"F��sz��Y�t���7�np�e�
%�hN��Z���3�/�ٓ�8��"��s}?H �歮�N�1[F3J�3_��5q�����,��0�/5
��P�5�t���7[�he�����ojZ"%`p�V^\�[hATZ��"���|i��8���3���S֣��/�Rpj�ܑ5g����tGj��uVlp38�FgX�%���?U���� �ݛ���Ѣ����F�PkdA�����܈W�N�k+�dl/<т�XD!�ёܝ�B���e�xַ��^SB���DV1�8��V?蓗4��L��2���k�F,�;n��u9�0;:]���]C4@sb����{�E��y7�]�3C�����CRb�▝�+3��X�V�>��sx��q{o�!͒=�K���t3�$LڴM]�"��7���N,m��@y�/��_!BS}S��1�lr��m.�[G�\���+\8�:�������� ��[-8VD �\b��.�vڙ�����K�8��?A��D�)�[���gC�Q �}���I�a�ӧw�ķ;�����%W�ki����*Ϛ����MV�&Hq1�8v��b�Α������-����`"GE�����{�b~���k�A�j��M=�@��YZl�}p'[Ul7z]�
yت*Cz�M=�;(�$�ݹF�S��~�!:�� �
{̠�f�Β�����!虇���c�3B�oyf���5K��w �ܽ�����]����A�5����o�*̨<PeNS�tI�F֬�RWND�P��
W֑�)�\�LL5��m��[�=X�ǕQG{��;Q��G�V��3m��;�暙Ԏ��Q���8��5����#h�O�B�	���A�RmuM��f�ޒa�+D�N���}�k�k^A��D������ʅ<vl���J������f��ދ��w8�Q��+5'���W��C; !���JZEXu5�`�[��<�u0g�r*�7Q�.��A�F+;!���tfF���W+�P!du@f33��T��w��E�Ay7)9*�À�>�apWC�;h�3u�#��
n�pG8N�0�4!�1�&i��;��W<�a��sX�a "�2+\LΉ,$�"j<Ӹ\	�8f���w���D�GO�j�Ƽ���z�I�J�͗&u
����eW�&nL�z�![`����1��[��T�Q��w�=?OQ��g�Y�&dT��!�s"ow��)5�(����>�-�l���9];86<����V?l�A��
�nj�MT- ��Q�Ywpp6
�uA̙���-��]�[z����+u���>,�獇p�P��G�Pa��M��,�wd��^����5t�	��#p����BG�}W�AhaM��#Kbf��jC���������ׇ�7"��o�U(�`��Zh�9������!�*
���$ ���~m�]%��*����S|_��z�Z�YP��_:&X���.���$+���P;56�8r�ne��d�� ������ Ӧ�[�"8/�7��.?-��C� K�Aբ�pY��t��H'R���D�HT��7�ȑ��̬�y�q�F�ޣ+���(֍zT6[��ƿj6#yvl:�e�c�y��U����VۚL��z3��$���i'v�G7�\L*��^�{���8�Nz>*���аegr��(��T>�F�Nj�}n�m�_��R3�=��]����Q� �u�^韼eև�Z!��\>Rզ���̌u�ΚR� ����~�����-i��@J�BE<�&��%\���?�C;��#ֻB��a��c���o��t��[��.�%���A�4��[��A�7~I����5Tj�Svff���G"7����*B�N
�8���������X~I�I`�w���fg/�6�M���m��4�JI知	}�a�?�p�\��:6�Ԋg�������Q��j��gIr�z ��r�:U�l������#{�B��2e�����%.���v�!�c
�zvg�O�yt��[VdŠ�N�A ı����N�dx���2Cr^��7P�d�
\�в���4�;`����:=��-ڡm;
���:.�f9�pw�##��Q�$���� `���ã!�QX�7���M�3�!�8hBSvS����"��ʻ��)��,bk��y�Q����D���e�&���ipy%��B����
@Ew��jf�����#���3�F����@I�Jǎ�*<\+�������YV(\G"O}�soC�I��㏖[1�	��aY$�����Y�ɔ��i���S�'� �õ$c���M�Z��$~�	Ԍ3��Oo�0|�@؛�PI�8�
��p��qK�ĜNO�0_������&�n�3�Ԫ}�-H�ɥ1���������Ɗ�h��p�	?��`I�ܩ��$�ez%> ��������-ִV�JĆ,�0��?��e�uH��\���5�pT�y�ҟ�4��D����ׅ��^�O��y�j���ٻ�~a:Sk��Y����IA^..@��2��@O� ׸�)�\1!y<%�[}z�u��kh�!�C�Q��*ٮӏS��s�c�S�9�Uf��;y��ˡ����ԟ`.�^9���<x�FH�mD�������X�w���h긤���g��Vb��Qmn60Q�q��k���&�C�]�~�Y\GtS��u��X�9�n�PQ��;�]^���d.u��^�ѕx���L�	�����ћM�ec�wf��[QU�U�z
/6���i�����q�hˌ5T��~ۃ���!1�RG�j�BI���L��S`��MD���������-���M'�A�O�:�]�o��2���X�TZ���a߷w�N�>FB�w��Y��=eg���� �����B��X=d6t.�n��[�#nd�6-�׏5I)9�cS�t�M%-ҐЂʉS��!N��^f!(Ѫ�8������,���X�%�>� �N�b�8�FNeYxw�=gi�hJj��5W�Vrg�Q�V��7�+e�Ku&1'^U$����`��@�Թx�j̚�g�����ua�f>�~c'�b������:M�,&�֞
Y:��V�7V�Qr�d�g�*�P�ϻ�]2���/�9��� 1�����1��t��q��}ZVPT�C������[�������Q�儜��(KV�����P��{b4i϶0�H��� =ε˩MfL+��m���?�(H���^���j�5fA�7\ W�mՓ'W�F�z9�{��	O�)��Rv��G����|��)�WV���0�EHa���3Q�q>(�rD�.5@%ᚲW�U?��Q�̉)�
�Ҫ�PT';�w�C	!,�t_��$P����l��3v<N��n8[��Ԁl��t?I���w�V�82���Yv7�~a$�A��!v�l,��	�ueAJ0�x�*|O������i�rp�|φ�by�t�7�z�_Q�l�R4t�"���'xC��C��$�Y@+۫Hk�dbwvdj⧜��~>� "���.�Iל,�>���b�Ƕ��2��W�eD�-���XK;�g�5��-�2}G�QZS�0S$w"N��n���h�λ}1C�qu9��Ǌ�u�[_ו��&z�Ҥx�� &�l���U��áѷ,���l���'�
TP�P�3����4�V;���_b�z��s�z�� $-��^$rcpÅ%�z��?fo�/(�נ��[L�#'R8�h"	�ҭ+~����V ��6@�4R	�KcՓu��%���{�`lB��8Ĭ@+�����8a�@���R�6���h��/������w[�_9�dw�3-Ih�l���7^J���\��h	�].��m:��r������bE�P$Ci`��ܻ�h�?�ƈ��ҥ��HV(V�nwkF�W�tn���R����*ۥ����R�-���H ������A��Ǉ���^�8����Ե��S���QK��@����見�sb��а��|y"V��N9�몃��h�'p%-��W[��W����3�L��=�'`c�$)����C�ڈ ���㈘�%>	U=�ң��X�eA�p�l7��Z�U��d->�O�j���O���E���?�����z��*ltd���N�xcd��|���DÆ�_m�E�݉z�����M�2����x����� (�Q:*SS9�n��TS�`�m#�dj�-� ݩ��>d{� ��?�,�<�`�_Ю����F ����U����}(�����+C�a�����*2�{������w!�bq�I�v�0�	X��ho��(
������=����~�\����kyh
y4��8��9�~<�,�:��$�5^,�/d��g?wD�f���� ���ۄ�(���Yݟx�W�t~���8�2>�B_r�1aJ��4OQ�<.[�H?'���s�W��ռ�ú�eR]JVD��Nr�m��:���qn��P�0k='�� ;m[��$m�1��(f�B�^���'���6]�׷��*�&��!�OD�n�́��n�5?�3��>�(���bu�d-AXb�X�s��m�(�U�?p�/.I�0g��N��c�w�2J���� R�Oବ�PAd��LM�n���47h�ކ�I�>R؜O5 ��~$z�y�qvփ��ڣ"�7�v�K;4o��vL<É�m��`�Լ�*#H��o\"�	 �8��x�n�;T@XF� 
�KVu�-��:R%����\]L8^�\�jv����SS� p�Zɓ���\���$C�zU��"�3ᕞG�7ñ��<@2]�t|c��`b���~�@A���%�op��)���W��8b�o����'�=�p-���)<1|X��5j�*-!�.��{9]+|�"�ͮ*f�m�D�u�hQ�FR���A� ����k�	�!��:	�x{Q�_���y�f���U�z��Ɨ���͗>Eg�,��H432{��վM)�
 A�f�x�Iu�l1w{/>�����,���;�����'@I@�P/���B�S���Nj��S�%1 ���6s�8�\�3���L�q�������������]�]=.&pY~�7p�Ź���P�%M7�}[Aq�ˈ�5��""C��	�HK�Э�Ǌ��*�7 ��������*wv�o���Z�	�d�7�J~{Ք���7�@��h��Q�]�v#�w��`��W���'�X%�tP�A�>�jY��mڌ#F o�]�P��O���2W�'
�n����i��E ݪO�i%���������I�#���)�+�F���>�+̍��F;}&:�ެ�#9 �6^0���;c�!
Lib!�y��д�'�,ږ��mvl��D��e��K�H*�{��_��޿3=����2f6P��nO����[͆/�?��r0���,;���TU�vs��{�~�6��훝�������{i-I$H�����l	ױ#MWb�T�X?�Y�4�8�U=ҺS��-��r�Ɲ)��U���L��ٿM-��&t)M:S��eL��!��U�"Ǆ�{��\Pɍ���̤�I�T��H5�0<��ٞsz���n'�T �DE\4�{E������^h�B���0n�6غ��!�Ie���>[���rΔ/k��	~��n���@�4�|v\�G��]yB�e�/���~����B�,�z:^;�D 2@5R�D�+ ��d�C,��n噑�b��޺>�0z:(�u��K=�����*T@�y)�̣l}s5�`�?�:���n�����Y����mGUK��eh�I�t���!�@����F���⑽��-�_�r��]��v5�8=���+bB��xv�Np��Ӑ�:�{��j)½��#�ʹvo�6�ݝ4��9 ��Dv����Մ�����$fz x �'13�S�V�Xc�ju��ۇ��*xÍK�)��rUC�=ֺ	c��Ud%�l1�a��)������ϡ�(J��▢7�]vᐻ7���U�M2;��9"{��kH��$�
ȇ���!c�ી�`����_�2ڥ|H�ݭ+�&�7Qa��>�7uV�/}���.����R+"��1��,��NJ�0	�.���d×�}��'ת11ʳo�"�le��xB�����?j�z���
y����o��p��֒4#4���5PV`��o��f���㭦�;O'�܆��՛�����<6�W<5bγF�ʌ;
�*3R�g��b��P�7����K���[���=�҆g�$#�(�V��߬ԋ����&��m�	���l�=�,����B,���]��C�]2��IƟ��n�@b`�e�c�i����Vz���7��:i��A.�|��a�ms7��[�9'r^�o����Dgom�ũ>r����y�a�{��g�g3������x�����)x�T����]j|R^ e2�,� [��£�q���]�覫�٤_�^ty}k�cf3oر*f��2D_}v�ա���b���pCc�(�"���p�(�Ju_��Z��,�NȐn$��6�j�C��"��QŸ��3�H`�����kP���f��J��O�﫰%�{�-e"p~j�u_7��D�&"S`[���u�	/&iA��g5�:!���j�b�#V79s>aLu�S��uoT?Ǻԟ�iH����m"@6�T|]��@?�C\��J*���_H�ڏ��僲 ����̦UE�3�y2�a8]Ð�����d�ٔ[��=���,6�6C������'^I��WUƁ(.t���\>�=��m9l�� �f�i�	Ѯ0�����������O��s&�=��z
,o���Һc-ө>��LM�%5L�Ue������^¥��StP[=5�\�_[�<���;U�d,��hL��Ϸf�e���9瘔�>M�r��6��
N��L�N^���u&,Pnʢ��.�C�q��,#�F�՘ɔT[m%�:��a�|%����˪G��"�C)��=XD�q�m���o��u��GFjY��!���vDGD�U�Nd��+�=eUiXkF=��6Z���O�1�a6R9�\���#l�O��Ǳ�0L����l��v�7q�